/*
    top.sv - Minimig on tang nano 20k toplevel
*/ 

/* we need two copies in case of 256k kickroms
     openFPGALoader --external-flash -o 0x400000 kick13.rom
     openFPGALoader --external-flash -o 0x440000 kick13.rom
   or a single copy of e.g. a 512k diag rom
     openFPGALoader --external-flash -o 0x400000 DiagROM
   or place a copy in the alternate rom slot (not supported yet)
     openFPGALoader --external-flash -o 0x480000 DiagROM   
*/
 
/* 
 TODO:
 - fix flash word counter
 - check why floppy sometimes hangs on boot
 - check why mouse counters sometimes go mad
 
 CHANGES:
 - remove userio
 - remove audio bitstream (sigma delta dac)
   - expose 14 bit digital interface (e.g. for HDMI)
 - remove ps2 keyboard from CIAA
   - expose CIAA keydat, keystrobe and keyack
   - bring keystrobe into 7Mhz clock domain
   - queue key events
   o (re-)implement caps lock
 - remove ps2 mouse from CIAA
   - expose digital mouse port
   - implement mouse event pointers
 - remove FPGA SPI from floppy.v
   - add generic sd card interface
   - expose sector interface to top
   - implement MFM encoding inside FPGA
  - remove sram_bridge
   - switch from ce to bank usage in sdram 
  
 */

module top(
  input			clk,

  input			reset, // button S2
  input			user,  // button S1

  output [5:0]	leds_n,
  output		ws2812,

  // spi flash interface
  output		mspi_cs,
  output		mspi_clk,
  inout			mspi_di,
  inout			mspi_hold,
  inout			mspi_wp,
  inout			mspi_do,

  // "Magic" port names that the gowin compiler connects to the on-chip SDRAM
  output		O_sdram_clk,
  output		O_sdram_cke,
  output		O_sdram_cs_n,  // chip select
  output		O_sdram_cas_n, // columns address select
  output		O_sdram_ras_n, // row address select
  output		O_sdram_wen_n, // write enable
  inout [31:0]	IO_sdram_dq, // 32 bit bidirectional data bus
  output [10:0]	O_sdram_addr, // 11 bit multiplexed address bus
  output [1:0]	O_sdram_ba, // two banks
  output [3:0]	O_sdram_dqm, // 32/4

  // generic IO, used for mouse/joystick/...
  input [7:0]	io,

  // interface to external BL616/M0S
  inout [5:0]	m0s,

  // MIDI/UART
  input			midi_in,
  output		midi_out,
		   
  // SD card slot
  output		sd_clk,
  inout			sd_cmd, // MOSI
  inout [3:0]	sd_dat, // 0: MISO
	   
  // SPI connection to ob-board BL616. By default an external
  // connection is used with a M0S Dock
  input			spi_sclk, // in... 
  input			spi_csn, // in (io?)
  output		spi_dir, // out
  input			spi_dat, // in (io?)

  // hdmi/tdms
  output		tmds_clk_n,
  output		tmds_clk_p,
  output [2:0]	tmds_d_n,
  output [2:0]	tmds_d_p
);

wire [5:0]	leds;
   
assign leds[5] = 1'b0;
assign leds_n = ~leds;  

// ============================== clock generation ===========================
   
// HDMI clock:  141.8758 MHz
// Pixel clock: 28.37516 MHz (HDMI/5)
// SDRAM clock: 70.9379 MHz (HDMI/2)
// Amiga clock: 7.09379 (Pixel/4)
   
`define PIXEL_CLOCK 28375160

wire clk_pixel_x5;   
wire pll_lock;   
pll_142m pll_hdmi (
    .clkout(clk_pixel_x5),
    .lock(pll_lock),
    .clkin(clk)
);

reg clk_71m;
always @(posedge clk_pixel_x5)
    clk_71m <= !clk_71m;

wire clk_pixel;
Gowin_CLKDIV clk_div_5 (
    .hclkin(clk_pixel_x5), // input hclkin
    .resetn(pll_lock),     // input resetn
    .clkout(clk_pixel)     // output clkout
);

wire	clk_28m = clk_pixel;

// generate 7 Mhz from 28Mhz
reg [1:0] clk_cnt;
always @(posedge clk_28m)
  clk_cnt <= clk_cnt + 2'd1;
   
wire	clk_7m = clk_cnt[1];

// control signals generated by the user via the OSD
wire 	osd_reset;   
   
// gemerate a reset for some time after rom has been initialized
reg [15:0] reset_cnt;
always @(posedge clk_7m) begin
    if(!rom_done || reset || osd_reset )
        reset_cnt <= 6'hffff;
    else if(reset_cnt != 0)
        reset_cnt = reset_cnt - 16'd1;
end

wire reset_i = |reset_cnt;
wire sdram_ready;

// -------------------------- M0S MCU interface -----------------------

// connect to ws2812 led
wire [23:0] ws2812_color;
ws2812 ws2812_inst (
    .clk(clk_28m),
    .color(ws2812_color),
    .data(ws2812)
);

// interface to M0S MCU
wire       mcu_sys_strobe;        // mcu message byte valid for sysctrl
wire       mcu_hid_strobe;        // -"- hid
wire       mcu_osd_strobe;        // -"- osd
wire       mcu_sdc_strobe;        // -"- sdc
wire       mcu_start;             // first byte of MCU message

wire [7:0] mcu_data_out;  

wire [7:0] sys_data_out;  
wire [7:0] hid_data_out;  
wire [7:0] osd_data_out = 8'h55;  // OSD actually has no data output
wire [7:0] sdc_data_out;

mcu_spi mcu (
	 .clk(clk_28m),
	 .reset(!pll_lock),

	 // SPI interface to BL616
     .spi_io_ss(m0s[2]),
     .spi_io_clk(m0s[3]),
     .spi_io_din(m0s[1]),
     .spi_io_dout(m0s[0]),

	 // byte wide data in/out to the submodules
     .mcu_sys_strobe(mcu_sys_strobe),
     .mcu_hid_strobe(mcu_hid_strobe),
     .mcu_osd_strobe(mcu_osd_strobe),
     .mcu_sdc_strobe(mcu_sdc_strobe),
     .mcu_start(mcu_start),
     .mcu_dout(mcu_data_out),
     .mcu_sys_din(sys_data_out),
     .mcu_hid_din(hid_data_out),
     .mcu_osd_din(osd_data_out),
     .mcu_sdc_din(sdc_data_out)
);

// decode SPI/MCU data received for human input devices (HID) and
// convert into Amiga compatible mouse and keyboard signals
wire [7:0] int_ack;
wire hid_int;
wire hid_iack = int_ack[1];
wire sdc_iack = int_ack[3];
wire [7:0] hid_joy0;   
   
// keyboard and mouse interface to Minimig
wire [5:0] mouse;  
wire       keystrobe;
wire [7:0] keydat;
wire       keyack;  

// signals to wire the floppy controller to the sd card
wire [3:0]  sd_rd;
wire [3:0]  sd_wr = 4'b0000;
wire [7:0]  sd_rd_data;
wire [7:0]  sd_wr_data = 8'h00;
wire [31:0] sd_sector;  
wire [8:0]  sd_byte_index;
wire        sd_rd_byte_strobe;
wire        sd_busy, sd_done;
wire [31:0] sd_img_size;
wire [3:0]  sd_img_mounted;
reg         sd_ready;
   
sd_card #(
    .CLK_DIV(3'd1)                   // for 28 Mhz clock
) sd_card (
    .rstn(pll_lock),                 // rstn active-low, 1:working, 0:reset
    .clk(clk_28m),                   // clock
  
    // SD card signals
    .sdclk(sd_clk),
    .sdcmd(sd_cmd),
    .sddat(sd_dat),

    // mcu interface
    .data_strobe(mcu_sdc_strobe),
    .data_start(mcu_start),
    .data_in(mcu_data_out),
    .data_out(sdc_data_out),

    // output file/image information. Image size is e.g. used by fdc to 
    // translate between sector/track/side and lba sector
    .image_mounted(sd_img_mounted),
    .image_size(sd_img_size),           // length of image file

    // interrupt to signal communication request
    .irq(sdc_int),
    .iack(sdc_iack),

    // user read sector command interface (sync with clk32)
    .rstart(sd_rd), 
    .wstart(sd_wr), 
    .rsector(sd_sector),
    .rbusy(sd_busy),
    .rdone(sd_done),

    // sector data output interface (sync with clk32)
    .inbyte(sd_wr_data),
    .outen(sd_rd_byte_strobe), // when outen=1, a byte of sector content is read out from outbyte
    .outaddr(sd_byte_index),   // outaddr from 0 to 511, because the sector size is 512
    .outbyte(sd_rd_data)       // a byte of sector content
);

hid hid (
        .clk(clk_28m),
        .reset(!pll_lock),

         // interface to receive user data from MCU (mouse, kbd, ...)
        .data_in_strobe(mcu_hid_strobe),
        .data_in_start(mcu_start),
        .data_in(mcu_data_out),
        .data_out(hid_data_out),

        // input local db9 port events to be sent to MCU. Changes also trigger
        // an interrupt, so the MCU doesn't have to poll for joystick events
        .db9_port( 6'h00 ),
        .irq( hid_int ),
        .iack( hid_iack ),

		.clk7(clk_7m),
        .mouse(mouse),
		 
        .keystrobe(keystrobe),
        .keydat(keydat),
        .keyack(keyack),
		 
        .joystick0(hid_joy0),
        .joystick1()
         );   

sysctrl sysctrl (
        .clk(clk_28m),
        .reset(!pll_lock),

         // interface to send and receive generic system control
        .data_in_strobe(mcu_sys_strobe),
        .data_in_start(mcu_start),
        .data_in(mcu_data_out),
        .data_out(sys_data_out),

        // values controlled by the OSD
        .system_reset(osd_reset),
        
        .int_out_n(m0s[4]),
        .int_in( { 4'b0000, sdc_int, 1'b0, hid_int, 1'b0 }),
        .int_ack( int_ack ),

        .buttons( {reset, user} ),
        .leds(),
        .color(ws2812_color)
);
   
// digital 12 bit video
wire hs_n, vs_n;
wire [3:0] red;
wire [3:0] green;
wire [3:0] blue;
   
wire [5:0] video_red;
wire [5:0] video_green;
wire [5:0] video_blue;   

osd_u8g2 osd_u8g2 (
        .clk(clk_28m),
        .reset(!pll_lock),

        .data_in_strobe(mcu_osd_strobe),
        .data_in_start(mcu_start),
        .data_in(mcu_data_out),

        .hs(hs_n),
        .vs(vs_n),
		     
        .r_in({red,   2'b00}),
        .g_in({green, 2'b00}),
        .b_in({blue,  2'b00}),
		     
        .r_out(video_red),
        .g_out(video_green),
        .b_out(video_blue)
);   

/* ---------------------- Minimig chipset ----------------------- */

// start cpu once the rom has been loaded from flash
wire    cpu_reset = !pll_lock || reset_i;

// two 15 bit audio channels
wire [14:0] audio_left;
wire [14:0] audio_right;   
  
// map first HID/USB joystick into second amiga joystick port
wire [5:0] n_joy2 = { !hid_joy0[5], !hid_joy0[4],
	  !hid_joy0[3], !hid_joy0[2], !hid_joy0[1], !hid_joy0[0] };   
   
wire [23:1] cpu_a;
wire cpu_as_n, cpu_lds_n, cpu_uds_n;
wire cpu_rw, cpu_dtack_n;
wire [2:0] ipl_n;
wire [15:0] cpu_din, cpu_dout;       

// Minimig ram/rom interface
wire [18:1] ram_a;
wire [15:0] ram_din;
wire [15:0] ram_dout;
wire [7:0]  ram_bank;    // 8 banks of 512k each
wire 	    ram_we_n;
wire [1:0]  ram_be;
wire 	    ram_oe_n;

wire [15:0] sdram_dout;

/* --------------------------- test rom/ram -------------------------- */

// using FPGA internal is useful if the external sdram/rom does not
// work reliably
   
// `define INTERNAL_MEM  // enable internal test memory (mainly rom)
// `define INTERNAL_RAM  // also enable so internal ram
   
`ifdef INTERNAL_MEM
reg [15:0] rom[0:1023];   // 2k rom
`ifdef INTERNAL_RAM
reg [15:0] ram[0:1023];   // 2k ram
`endif   
initial begin
    $readmemh ("ram_test/ram_test.hex", rom, 0);
end

// memory io stats oen cycle after start of 7mhz rising edge
reg [15:0] mem_dout;
always @(posedge clk_28m)
    mem_dout <= 
        (ram_bank[3])?rom[ram_a[10:1]]:
`ifdef INTERNAL_RAM
        (ram_bank[0])?ram[ram_a[10:1]]:
`endif
        16'h0000;

`ifdef INTERNAL_RAM
// ram write happens in the middle of the 7Mhz cycle
always @(negedge clk_7m)
    if(ram_bank[0] && !ram_we_n && ram_a[18:11]==8'h00)
        ram[ram_a[10:1]] <= ram_dout;

// with internal ram _all_ memory access in the first 2k go internal
wire	   mem_access = ram_a[18:11]==8'h00;  
`else
// without internal ram only the first 2k ROM access is internal
wire	   mem_access = ram_bank[3] && ram_a[18:11]==8'h00;     
`endif

// map internal memory to first 2k of kickstart/chipram space
// address lines 18:1 are valid with each 512k block
assign ram_din = mem_access?mem_dout:sdram_dout;
`else
assign ram_din = sdram_dout;
`endif

Minimig1 MINIMIG1 
(
   // m68k pins
   .cpu_address(cpu_a),       // m68k address bus
   .cpu_data(cpu_din),        // m68k data bus
   .cpu_wrdata(cpu_dout),     // m68k data bus
   .n_cpu_ipl(ipl_n),         // m68k interrupt request
   .n_cpu_as(cpu_as_n),       // m68k address strobe
   .n_cpu_uds(cpu_uds_n),     // m68k upper data strobe
   .n_cpu_lds(cpu_lds_n),     // m68k lower data strobe
   .cpu_r_w(cpu_rw),          // m68k read / write
   .n_cpu_dtack(cpu_dtack_n), // m68k data acknowledge
   
   // sram pins
   .ram_data(ram_dout),       // sram data bus
   .ram_address_out(ram_a),   // sram address bus
   .ramdata_in(ram_din),      // sram data bus in
   .bank(ram_bank),           // ram/rom bank
   .n_ram_bhe(ram_be[1]),     // sram upper byte select
   .n_ram_ble(ram_be[0]),     // sram lower byte select
   .n_ram_we(ram_we_n),       // sram write enable
   .n_ram_oe(ram_oe_n),       // sram output enable
   
   // system pins
   .clk(clk_7m),      // system clock (7.09379 MHz)
   .clk28m(clk_28m),  // 28.37516 MHz clock

   // rs232 pins are connected to the pins used for MIDI on Atari ST
   // connecting a USB UART adapter here allows to e.g. control DiagROM from a PC
   .rxd(midi_in),     // rs232 receive
   .txd(midi_out),    // rs232 send
   .cts(1'b1),        // rs232 clear to send
   .rts(),            // rs232 request to send
   
   // I/O
   .n_joy1(6'h3f),     // joystick 1 [fire2,fire,right,left,down,up] (default mouse port)
   .n_joy2(n_joy2),    // joystick 2 [fire2,fire,right,left,down,up] (default joystick port)
   .n_15khz(1'b1),     // scandoubler is permanently enabled
   .pwrled(leds[0]),   // power led

   // keyboard and mouse event input
   .keystrobe(keystrobe),
   .keydat(keydat),
   .keyack(keyack),
   .mouse(mouse),
 
   // video
   .n_hsync(hs_n),     // horizontal sync
   .n_vsync(vs_n),     // vertical sync
   .red(red),          // red
   .green(green),      // green
   .blue(blue),        // blue
   
   // audio
   .aud_l(audio_left),   // left DAC data
   .aud_r(audio_right),  // right DAC data
 
    // sd card interface for floppy disk emulation
   .sdc_img_size(sd_img_size),
   .sdc_img_mounted(sd_img_mounted), 
   .sdc_rd(sd_rd),
   .sdc_sector(sd_sector),
   .sdc_busy(sd_busy),
   .sdc_done(sd_done), 
   .sdc_byte_in_strobe(sd_rd_byte_strobe),
   .sdc_byte_in_addr(sd_byte_index),
   .sdc_byte_in_data(sd_rd_data),
  
   // user i/o
   .floppyled(leds[1]),
   
   // unused pins
   .cpurst(cpu_reset),
   .n_joy3(5'h1f),      // joystick 3 [fire2,fire,right,left,down,up] (printer port)
   .n_joy4(5'h1f)       // joystick 4 [fire2,fire,right,left,down,up] (printer port)
);

/* ------------------- fx68k cycle exact CPU core  ------------------- */
reg  phi1, phi2;   
   
always @(posedge clk_28m) begin
   if(cpu_reset) begin
	  phi1 <= 0;
	  phi2 <= 0;
   end else begin   
	  phi1 <= 0;
	  phi2 <= 0;
	  if(clk_cnt[0] &&  clk_cnt[1]) phi1 <= 1;   
	  if(clk_cnt[0] && ~clk_cnt[1]) phi2 <= 1;
   end
end

fx68k fx68k (
     .clk        ( clk_28m     ),
     .extReset   ( cpu_reset   ),
     .pwrUp      ( reset       ),
     .enPhi1     ( phi1        ),
     .enPhi2     ( phi2        ),
     .eRWn       ( cpu_rw      ),
     .ASn        ( cpu_as_n    ),
     .LDSn       ( cpu_lds_n   ),
     .UDSn       ( cpu_uds_n   ),
     .E          (             ),
     .VMAn       (             ),
     .FC0        (             ),
     .FC1        (             ),
     .FC2        (             ),
     .BGn        (             ),
     .oRESETn    (             ),
     .oHALTEDn   (             ),
     .DTACKn     ( cpu_dtack_n ),
     .VPAn       ( 1'b1        ),
     .BERRn      ( 1'b1        ),
     .HALTn      ( 1'b1        ),
     .BRn        ( 1'b1        ),
     .BGACKn     ( 1'b1        ),
     .IPL0n      ( ipl_n[0]    ),
     .IPL1n      ( ipl_n[1]    ),
     .IPL2n      ( ipl_n[2]    ),
     .iEdb       ( cpu_din     ),
     .oEdb       ( cpu_dout    ),
     .eab        ( cpu_a       )
);

wire           flash_ready;  
wire           mem_ready = sdram_ready && flash_ready && pll_lock;  
   
reg            start_rom_copy;
reg            mem_ready_D;

// geneate a start_rom_copy signal once flash and SDRAM are initialized
always @(posedge clk_28m or negedge pll_lock) begin
   if(!pll_lock) begin
      start_rom_copy <= 1'b0;
      mem_ready_D <= 1'b0;
         
   end else begin
      mem_ready_D <= mem_ready;  
      start_rom_copy <= 1'b0;         

      if(mem_ready && !mem_ready_D)
          start_rom_copy <= 1'b1;     
   end
end

/* -------------- state machine copying data from flash to sdram ---------------- */
reg [21:0]  flash_addr;  
wire [15:0] flash_dout;
reg [15:0]  flash_doutD;
reg		    flash_cs;  
reg [31:0]  word_count;
reg [2:0]   state;
wire        flash_data_strobe;
wire        flash_busy;   

// once the copy counter has run to zero, all rom has been copied
wire		rom_done = (word_count == 0);

assign leds[4] = !pll_lock;   
assign leds[3] = !mem_ready;  
assign leds[2] = !rom_done;  
   
reg [21:0]  flash_ram_addr;   
reg         flash_ram_write;
reg [5:0]   flash_cnt;  

always @(posedge clk_28m or negedge mem_ready) begin
    if(!mem_ready) begin
       flash_addr <= 22'h200000;          // 4MB flash offset (word address)
       flash_ram_addr <= { 4'h1, 18'h0 }; // write into 512k sdram segment used for kick rom
       word_count <= 22'h40001;           // 512k bytes ROM data = 256k words

       state <= 3'h0;
       flash_ram_write <= 1'b0;
       flash_cs <= 1'b0;        
       flash_cnt <= 6'd0;
    end else begin
        if((start_rom_copy || state == 7) && (word_count != 0)) begin
            flash_cs <= 1'b1;
            flash_cnt <= 6'd15; // >= 30 @ 32MHz
        end else begin
            if(flash_cnt != 0) flash_cnt <= flash_cnt - 6'd1;
            if(flash_busy)     flash_cs <= 1'b0;

            // ... static timing with fixed counter
            if(flash_cnt == 6'd1) begin
                state <= 1;
                flash_addr <= flash_addr + 22'd1;
                word_count <= word_count - 22'd1;

                // we don't necessarily need to latch the data. But latching it here
                // allows to exactly determine the real access time by adjusting flash_cnt
                // to the lowest value that gives a stable image
                flash_doutD <= flash_dout;
            end
        end

        // advance ram write state
        if(state != 0)  state <= state + 3'd1;
        if(state == 1)  flash_ram_write <= 1'b1;
        if(state == 6)  flash_ram_write <= 1'b0;
        if(state == 7)  flash_ram_addr <= flash_ram_addr + 22'd1;
    end
end

// ----------------------------- SDRAM ---------------------------------

assign O_sdram_addr = sd_addr[10:0];
wire [12:0] sd_addr;

// sdram can be addressed during runtime by minimig and at startup
// by flash rom loader

// RAM banks are:
// 0 - 0000 0001 - chip0
// 1 - 0000 0010 - chip1
// 2 - 0000 0100 - chip2
// 3 - 0000 1000 - kick
// 4 - 0001 0000 - slow0
// 5 - 0010 0000 - chip3
// 6 - 0100 0000 - slow2
// 7 - 1000 0000 - slow1
   
// there's a total of 16 sdram segments of 512kBytes
// enable sdram for up to 2MB chip and 512k kick
wire [3:0] sdram_segment = 
		   (ram_bank == 8'b0000_0001)?4'h0:    // chip0
		   (ram_bank == 8'b0000_1000)?4'h1:    // kick
		   (ram_bank == 8'b0000_0010)?4'h2:    // chip1
		   (ram_bank == 8'b0000_0100)?4'h3:    // chip2
		   (ram_bank == 8'b0010_0000)?4'h4:    // chip3
		   (ram_bank == 8'b0001_0000)?4'h5:    // slow0
		   (ram_bank == 8'b1000_0000)?4'h6:    // slow1
		   (ram_bank == 8'b0100_0000)?4'h7:    // slow2
		   4'hf;

wire    sdram_access = ram_bank != 0;  
wire    sdram_rw     = sdram_access && (ram_bank != 8) && !ram_we_n;  

wire		sdram_refresh = rom_done?!sdram_access:1'b0;
wire [21:0] sdram_addr    = rom_done?{sdram_segment,ram_a}:flash_ram_addr;
wire [15:0] sdram_din     = rom_done?ram_dout:flash_doutD;
wire [1:0]  sdram_be      = rom_done?ram_be:2'b00;
wire		sdram_cs      = rom_done?clk_7m:flash_ram_write;
wire		sdram_we      = rom_done?sdram_rw:flash_ram_write; 
   
sdram sdram (
  	.sd_clk     ( O_sdram_clk   ), // sd clock
	.sd_cke     ( O_sdram_cke   ), // clock enable
	.sd_data    ( IO_sdram_dq   ), // 32 bit bidirectional data bus
	.sd_addr    ( sd_addr       ), // 11 bit multiplexed address bus
	.sd_dqm     ( O_sdram_dqm   ), // two byte masks
	.sd_ba      ( O_sdram_ba    ), // two banks
	.sd_cs      ( O_sdram_cs_n  ), // a single chip select
	.sd_we      ( O_sdram_wen_n ), // write enable
	.sd_ras     ( O_sdram_ras_n ), // row address select
	.sd_cas     ( O_sdram_cas_n ), // columns address select

	// cpu/chipset interface
	.clk        ( clk_71m       ), // sdram is accessed at 71MHz
	.reset_n    ( pll_lock      ), // init signal after FPGA config to initialize RAM

	.ready      ( sdram_ready   ), // ram is ready and has been initialized
	.refresh    ( sdram_refresh ), // chipset requests a refresh cycle
	.din        ( sdram_din     ), // data input from chipset/cpu
	.dout       ( sdram_dout    ),
	.addr       ( sdram_addr    ), // 22 bit word address
	.ds         ( sdram_be      ), // upper/lower data strobe
	.cs         ( sdram_cs      ), // cpu/chipset requests read/wrie
	.we         ( sdram_we      )  // cpu/chipset requests write
);

// run the flash a 71MHz. This is only used at power-up to copy kickstart
// from flash to sdram
assign mspi_clk = ~clk_71m;   
flash flash (
    .clk       ( clk_71m     ),
    .resetn    ( pll_lock    ),
    .ready     ( flash_ready ),

    .address   ( flash_addr  ),
    .cs        ( flash_cs    ),
    .dout      ( flash_dout  ),
	.busy      ( flash_busy  ),

    .mspi_cs   ( mspi_cs     ),
    .mspi_di   ( mspi_di     ),
    .mspi_hold ( mspi_hold   ),
    .mspi_wp   ( mspi_wp     ),
    .mspi_do   ( mspi_do     )
);

/* -------------------- HDMI video and audio -------------------- */

// generate 48khz audio clock
reg clk_audio;
reg [8:0] aclk_cnt;
always @(posedge clk_pixel) begin
    // divisor = pixel clock / 48000 / 2 - 1
    if(aclk_cnt < `PIXEL_CLOCK / 48000 / 2 -1)
        aclk_cnt <= aclk_cnt + 9'd1;
    else begin
        aclk_cnt <= 9'd0;
        clk_audio <= ~clk_audio;
    end
end
   
wire [2:0] tmds;
wire tmds_clock;

wire vreset;
video_analyzer video_analyzer (
    .clk    ( clk_28m ),
    .hs     ( hs_n    ),
    .vs     ( vs_n    ),
    .vreset ( vreset  )
);
   
hdmi #(
    .AUDIO_RATE(48000), .AUDIO_BIT_WIDTH(16),
    .VENDOR_NAME( { "MiSTle", 16'd0} ),
    .PRODUCT_DESCRIPTION( {"Nanomig", 72'd0} )
) hdmi(
  .clk_pixel_x5(clk_pixel_x5),
  .clk_pixel(clk_pixel),
  .clk_audio(clk_audio),
  .audio_sample_word( { { 1'b0, ~audio_left[14],audio_left[13:0]}, {1'b0, ~audio_right[14],audio_right[13:0]}} ),
  .tmds(tmds),
  .tmds_clock(tmds_clock),

  .reset(vreset),    // signal to synchronize HDMI

  .rgb( { video_red, 2'b00, video_green, 2'b00, video_blue, 2'b00 } )
);

// differential output
ELVDS_OBUF tmds_bufds [3:0] (
        .I({tmds_clock, tmds}),
        .O({tmds_clk_p, tmds_d_p}),
        .OB({tmds_clk_n, tmds_d_n})
);
   
endmodule

// To match emacs with gw_ide default
// Local Variables:
// tab-width: 4
// End:

