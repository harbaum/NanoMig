module tg68k_alu_2_1_2_1
  (input  clk,
   input  reset,
   input  clkena_lw,
   input  [1:0] cpu,
   input  execopc,
   input  decodeopc,
   input  exe_condition,
   input  exec_tas,
   input  long_start,
   input  non_aligned,
   input  check_aligned,
   input  movem_presub,
   input  set_stop,
   input  z_error,
   input  [1:0] rot_bits,
   input  [88:0] exec,
   input  [31:0] op1out,
   input  [31:0] op2out,
   input  [31:0] reg_qa,
   input  [31:0] reg_qb,
   input  [15:0] opcode,
   input  [15:0] exe_opcode,
   input  [1:0] exe_datatype,
   input  [15:0] sndopc,
   input  [15:0] last_data_read,
   input  [15:0] data_read,
   input  [7:0] flagssr,
   input  [6:0] micro_state,
   input  [7:0] bf_ext_in,
   input  [5:0] bf_shift,
   input  [5:0] bf_width,
   input  [31:0] bf_ffo_offset,
   input  [4:0] bf_loffset,
   output [7:0] bf_ext_out,
   output set_v_flag,
   output [7:0] flags,
   output [2:0] c_out,
   output [31:0] addsub_q,
   output [31:0] aluout);
  wire [31:0] op1in;
  wire [31:0] addsub_a;
  wire [31:0] addsub_b;
  wire [33:0] notaddsub_b;
  wire [33:0] add_result;
  wire [2:0] addsub_ofl;
  wire opaddsub;
  wire [3:0] c_in;
  wire [2:0] flag_z;
  wire [3:0] set_flags;
  wire [7:0] ccrin;
  wire [3:0] last_flags1;
  wire [9:0] bcd_pur;
  wire [8:0] bcd_kor;
  wire halve_carry;
  wire vflag_a;
  wire bcd_a_carry;
  wire [8:0] bcd_a;
  wire [127:0] result_mulu;
  wire [63:0] result_div;
  wire [31:0] result_div_pre;
  wire set_mv_flag;
  wire v_flag;
  wire rot_rot;
  wire rot_x;
  wire rot_c;
  wire [31:0] rot_out;
  wire asl_vflag;
  wire [4:0] bit_number;
  wire [31:0] bits_out;
  wire one_bit_in;
  wire bchg;
  wire bset;
  wire [63:0] mulu_reg;
  wire [31:0] faktora;
  wire [31:0] faktorb;
  wire [63:0] div_reg;
  wire [63:0] div_quot;
  wire div_neg;
  wire div_bit;
  wire [32:0] div_sub;
  wire [32:0] div_over;
  wire nozero;
  wire div_qsign;
  wire [63:0] dividend;
  wire divs;
  wire signedop;
  wire op1_sign;
  wire [15:0] op2outext;
  wire [31:0] datareg;
  wire [31:0] bf_datareg;
  wire [39:0] result;
  wire [39:0] result_tmp;
  wire [31:0] unshifted_bitmask;
  wire [39:0] inmux0;
  wire [39:0] inmux1;
  wire [39:0] inmux2;
  wire [31:0] inmux3;
  wire [39:0] shifted_bitmask;
  wire [37:0] bitmaskmux0;
  wire [35:0] bitmaskmux1;
  wire [31:0] bitmaskmux2;
  wire [31:0] bitmaskmux3;
  wire [31:0] bf_set2;
  wire [39:0] shift;
  wire [5:0] bf_firstbit;
  wire [3:0] mux;
  wire [4:0] bitnr;
  wire [31:0] mask;
  wire mask_not_zero;
  wire bf_bset;
  wire bf_nflag;
  wire bf_bchg;
  wire bf_ins;
  wire bf_exts;
  wire bf_fffo;
  wire bf_d32;
  wire bf_s32;
  wire [33:0] hot_msb;
  wire [32:0] vector;
  wire [65:0] result_bs;
  wire [5:0] bit_nr;
  wire [5:0] bit_msb;
  wire [5:0] bs_shift;
  wire [5:0] bs_shift_mod;
  wire [32:0] asl_over;
  wire [32:0] asl_over_xor;
  wire [32:0] asr_sign;
  wire msb;
  wire [5:0] ring;
  wire [31:0] alu;
  wire [31:0] bsout;
  wire bs_v;
  wire bs_c;
  wire bs_x;
  wire n9536_o;
  wire n9537_o;
  wire [23:0] n9538_o;
  wire [6:0] n9539_o;
  wire n9540_o;
  wire [31:0] n9541_o;
  wire [31:0] n9542_o;
  wire [31:0] n9543_o;
  wire [31:0] n9544_o;
  wire [31:0] n9545_o;
  wire [31:0] n9546_o;
  wire n9547_o;
  wire n9548_o;
  wire n9549_o;
  wire [7:0] n9550_o;
  wire n9551_o;
  wire n9553_o;
  wire n9554_o;
  wire [31:0] n9555_o;
  wire [31:0] n9556_o;
  wire [31:0] n9557_o;
  wire n9558_o;
  wire n9560_o;
  wire n9561_o;
  wire n9563_o;
  wire [15:0] n9564_o;
  wire [15:0] n9565_o;
  wire [31:0] n9566_o;
  wire n9567_o;
  wire [31:0] n9568_o;
  wire [31:0] n9569_o;
  wire [31:0] n9570_o;
  wire [31:0] n9571_o;
  wire n9572_o;
  wire [31:0] n9573_o;
  wire n9574_o;
  wire [31:0] n9575_o;
  wire n9576_o;
  wire [3:0] n9577_o;
  wire [3:0] n9578_o;
  wire [7:0] n9579_o;
  wire n9580_o;
  wire [31:0] n9581_o;
  wire n9582_o;
  wire n9583_o;
  wire n9584_o;
  wire n9585_o;
  wire [15:0] n9586_o;
  wire [15:0] n9587_o;
  wire [31:0] n9588_o;
  wire n9589_o;
  wire n9590_o;
  wire n9591_o;
  wire n9592_o;
  wire [7:0] n9594_o;
  wire n9595_o;
  wire [3:0] n9596_o;
  wire [3:0] n9597_o;
  wire [7:0] n9598_o;
  wire [7:0] n9599_o;
  wire [7:0] n9600_o;
  wire [15:0] n9601_o;
  wire [7:0] n9602_o;
  wire [7:0] n9603_o;
  wire [7:0] n9604_o;
  wire [7:0] n9605_o;
  wire [7:0] n9606_o;
  wire [15:0] n9607_o;
  wire [15:0] n9608_o;
  wire [15:0] n9609_o;
  wire [15:0] n9610_o;
  wire [15:0] n9611_o;
  wire [15:0] n9612_o;
  wire [31:0] n9613_o;
  wire [31:0] n9614_o;
  wire [31:0] n9615_o;
  wire [31:0] n9616_o;
  wire [31:0] n9617_o;
  wire [31:0] n9618_o;
  wire [31:0] n9619_o;
  wire [7:0] n9620_o;
  wire [7:0] n9621_o;
  wire [23:0] n9622_o;
  wire [23:0] n9623_o;
  wire [23:0] n9624_o;
  wire [31:0] n9625_o;
  wire [31:0] n9626_o;
  wire [31:0] n9627_o;
  wire [31:0] n9628_o;
  wire [31:0] n9629_o;
  wire [7:0] n9630_o;
  wire [7:0] n9631_o;
  wire [23:0] n9632_o;
  wire [23:0] n9633_o;
  wire [23:0] n9634_o;
  wire n9639_o;
  wire n9640_o;
  wire n9641_o;
  wire n9642_o;
  wire [1:0] n9643_o;
  wire n9644_o;
  wire [2:0] n9645_o;
  wire [28:0] n9646_o;
  wire [31:0] n9647_o;
  wire [1:0] n9648_o;
  wire [31:0] n9650_o;
  wire [31:0] n9651_o;
  wire [31:0] n9652_o;
  wire n9653_o;
  wire n9656_o;
  wire n9658_o;
  wire [3:0] n9659_o;
  wire [7:0] n9661_o;
  wire [11:0] n9663_o;
  wire [3:0] n9664_o;
  wire [15:0] n9665_o;
  wire n9666_o;
  wire n9667_o;
  wire n9668_o;
  wire n9669_o;
  wire n9670_o;
  wire n9671_o;
  wire n9672_o;
  wire n9673_o;
  wire n9675_o;
  wire n9676_o;
  wire n9677_o;
  wire n9678_o;
  wire n9679_o;
  wire n9680_o;
  wire n9682_o;
  wire n9683_o;
  wire n9684_o;
  wire n9685_o;
  wire n9686_o;
  wire n9687_o;
  wire n9688_o;
  wire n9689_o;
  wire [31:0] n9692_o;
  wire [31:0] n9694_o;
  wire [31:0] n9696_o;
  wire n9697_o;
  wire n9698_o;
  wire n9699_o;
  wire n9700_o;
  wire n9701_o;
  wire n9703_o;
  wire n9704_o;
  wire [31:0] n9705_o;
  wire n9706_o;
  wire n9707_o;
  wire [15:0] n9708_o;
  wire [15:0] n9709_o;
  wire [15:0] n9710_o;
  wire [15:0] n9711_o;
  wire [15:0] n9712_o;
  wire n9714_o;
  wire n9715_o;
  wire n9716_o;
  wire n9717_o;
  wire n9718_o;
  wire n9719_o;
  wire n9720_o;
  wire [31:0] n9722_o;
  wire [31:0] n9723_o;
  wire n9724_o;
  wire n9725_o;
  wire n9727_o;
  wire [31:0] n9730_o;
  wire [31:0] n9731_o;
  wire [31:0] n9732_o;
  wire [31:0] n9733_o;
  wire [31:0] n9734_o;
  wire [31:0] n9735_o;
  wire n9736_o;
  wire n9737_o;
  wire [32:0] n9739_o;
  wire n9740_o;
  wire [33:0] n9741_o;
  wire [32:0] n9743_o;
  wire n9744_o;
  wire [33:0] n9745_o;
  wire [33:0] n9746_o;
  wire [33:0] n9747_o;
  wire [32:0] n9749_o;
  wire n9750_o;
  wire [33:0] n9751_o;
  wire [33:0] n9752_o;
  wire n9753_o;
  wire n9754_o;
  wire n9755_o;
  wire n9756_o;
  wire n9757_o;
  wire n9758_o;
  wire n9759_o;
  wire n9760_o;
  wire n9761_o;
  wire n9762_o;
  wire n9763_o;
  wire [31:0] n9764_o;
  wire n9765_o;
  wire n9766_o;
  wire n9767_o;
  wire n9768_o;
  wire n9769_o;
  wire n9770_o;
  wire n9771_o;
  wire n9772_o;
  wire n9773_o;
  wire n9774_o;
  wire n9775_o;
  wire n9776_o;
  wire n9777_o;
  wire n9778_o;
  wire n9779_o;
  wire n9780_o;
  wire n9781_o;
  wire n9782_o;
  wire n9783_o;
  wire n9784_o;
  wire n9785_o;
  wire [2:0] n9786_o;
  wire n9790_o;
  wire [8:0] n9791_o;
  wire [9:0] n9792_o;
  wire n9793_o;
  wire n9794_o;
  wire n9795_o;
  wire n9796_o;
  wire n9797_o;
  wire [3:0] n9800_o;
  localparam [8:0] n9801_o = 9'b000000000;
  wire n9803_o;
  wire [3:0] n9805_o;
  wire [3:0] n9806_o;
  wire n9807_o;
  wire n9808_o;
  wire n9809_o;
  wire n9810_o;
  wire n9811_o;
  wire n9812_o;
  wire [8:0] n9813_o;
  wire [8:0] n9814_o;
  wire n9815_o;
  wire n9816_o;
  wire n9817_o;
  wire n9818_o;
  wire n9819_o;
  wire [3:0] n9821_o;
  wire n9822_o;
  wire n9823_o;
  wire n9824_o;
  wire n9825_o;
  wire n9826_o;
  wire n9827_o;
  wire n9828_o;
  wire n9829_o;
  wire n9830_o;
  wire n9831_o;
  wire n9832_o;
  wire n9833_o;
  wire n9834_o;
  wire [3:0] n9836_o;
  wire n9837_o;
  wire n9838_o;
  wire n9839_o;
  wire n9840_o;
  wire [8:0] n9841_o;
  wire [8:0] n9842_o;
  wire [7:0] n9843_o;
  wire [7:0] n9844_o;
  wire [7:0] n9845_o;
  wire n9846_o;
  wire [8:0] n9847_o;
  wire n9848_o;
  wire n9850_o;
  wire n9851_o;
  wire n9852_o;
  wire n9853_o;
  wire [1:0] n9858_o;
  wire n9860_o;
  wire n9862_o;
  wire [1:0] n9863_o;
  reg n9866_o;
  reg n9870_o;
  wire n9876_o;
  wire n9877_o;
  wire [1:0] n9878_o;
  wire n9880_o;
  wire [4:0] n9881_o;
  wire [2:0] n9882_o;
  wire [4:0] n9884_o;
  wire [4:0] n9885_o;
  wire [1:0] n9886_o;
  wire n9888_o;
  wire [4:0] n9889_o;
  wire [2:0] n9890_o;
  wire [4:0] n9892_o;
  wire [4:0] n9893_o;
  wire [4:0] n9894_o;
  wire n9900_o;
  wire n9901_o;
  wire n9902_o;
  wire [1:0] n9908_o;
  wire n9910_o;
  wire n9913_o;
  wire [2:0] n9915_o;
  wire n9917_o;
  wire n9919_o;
  wire n9921_o;
  wire n9923_o;
  wire n9925_o;
  wire [4:0] n9926_o;
  reg n9929_o;
  reg n9933_o;
  reg n9937_o;
  reg n9941_o;
  reg n9945_o;
  reg n9948_o;
  wire [1:0] n9949_o;
  wire n9951_o;
  wire n9954_o;
  wire [7:0] n9956_o;
  wire [4:0] n9974_o;
  wire n9976_o;
  wire n9979_o;
  wire n9980_o;
  wire n9981_o;
  wire n9982_o;
  wire n9987_o;
  localparam [31:0] n9988_o = 32'b00000000000000000000000000000000;
  wire [4:0] n9990_o;
  wire n9992_o;
  wire n9995_o;
  wire n9996_o;
  wire n9997_o;
  wire n9998_o;
  wire n10002_o;
  wire n10003_o;
  wire [4:0] n10005_o;
  wire n10007_o;
  wire n10010_o;
  wire n10011_o;
  wire n10012_o;
  wire n10013_o;
  wire n10017_o;
  wire n10018_o;
  wire [4:0] n10020_o;
  wire n10022_o;
  wire n10025_o;
  wire n10026_o;
  wire n10027_o;
  wire n10028_o;
  wire n10032_o;
  wire n10033_o;
  wire [4:0] n10035_o;
  wire n10037_o;
  wire n10040_o;
  wire n10041_o;
  wire n10042_o;
  wire n10043_o;
  wire n10047_o;
  wire n10048_o;
  wire [4:0] n10050_o;
  wire n10052_o;
  wire n10055_o;
  wire n10056_o;
  wire n10057_o;
  wire n10058_o;
  wire n10062_o;
  wire n10063_o;
  wire [4:0] n10065_o;
  wire n10067_o;
  wire n10070_o;
  wire n10071_o;
  wire n10072_o;
  wire n10073_o;
  wire n10077_o;
  wire n10078_o;
  wire [4:0] n10080_o;
  wire n10082_o;
  wire n10085_o;
  wire n10086_o;
  wire n10087_o;
  wire n10088_o;
  wire n10092_o;
  wire n10093_o;
  wire [4:0] n10095_o;
  wire n10097_o;
  wire n10100_o;
  wire n10101_o;
  wire n10102_o;
  wire n10103_o;
  wire n10107_o;
  wire n10108_o;
  wire [4:0] n10110_o;
  wire n10112_o;
  wire n10115_o;
  wire n10116_o;
  wire n10117_o;
  wire n10118_o;
  wire n10122_o;
  wire n10123_o;
  wire [4:0] n10125_o;
  wire n10127_o;
  wire n10130_o;
  wire n10131_o;
  wire n10132_o;
  wire n10133_o;
  wire n10137_o;
  wire n10138_o;
  wire [4:0] n10140_o;
  wire n10142_o;
  wire n10145_o;
  wire n10146_o;
  wire n10147_o;
  wire n10148_o;
  wire n10152_o;
  wire n10153_o;
  wire [4:0] n10155_o;
  wire n10157_o;
  wire n10160_o;
  wire n10161_o;
  wire n10162_o;
  wire n10163_o;
  wire n10167_o;
  wire n10168_o;
  wire [4:0] n10170_o;
  wire n10172_o;
  wire n10175_o;
  wire n10176_o;
  wire n10177_o;
  wire n10178_o;
  wire n10182_o;
  wire n10183_o;
  wire [4:0] n10185_o;
  wire n10187_o;
  wire n10190_o;
  wire n10191_o;
  wire n10192_o;
  wire n10193_o;
  wire n10197_o;
  wire n10198_o;
  wire [4:0] n10200_o;
  wire n10202_o;
  wire n10205_o;
  wire n10206_o;
  wire n10207_o;
  wire n10208_o;
  wire n10212_o;
  wire n10213_o;
  wire [4:0] n10215_o;
  wire n10217_o;
  wire n10220_o;
  wire n10221_o;
  wire n10222_o;
  wire n10223_o;
  wire n10227_o;
  wire n10228_o;
  wire [4:0] n10230_o;
  wire n10232_o;
  wire n10235_o;
  wire n10236_o;
  wire n10237_o;
  wire n10238_o;
  wire n10242_o;
  wire n10243_o;
  wire [4:0] n10245_o;
  wire n10247_o;
  wire n10250_o;
  wire n10251_o;
  wire n10252_o;
  wire n10253_o;
  wire n10257_o;
  wire n10258_o;
  wire [4:0] n10260_o;
  wire n10262_o;
  wire n10265_o;
  wire n10266_o;
  wire n10267_o;
  wire n10268_o;
  wire n10272_o;
  wire n10273_o;
  wire [4:0] n10275_o;
  wire n10277_o;
  wire n10280_o;
  wire n10281_o;
  wire n10282_o;
  wire n10283_o;
  wire n10287_o;
  wire n10288_o;
  wire [4:0] n10290_o;
  wire n10292_o;
  wire n10295_o;
  wire n10296_o;
  wire n10297_o;
  wire n10298_o;
  wire n10302_o;
  wire n10303_o;
  wire [4:0] n10305_o;
  wire n10307_o;
  wire n10310_o;
  wire n10311_o;
  wire n10312_o;
  wire n10313_o;
  wire n10317_o;
  wire n10318_o;
  wire [4:0] n10320_o;
  wire n10322_o;
  wire n10325_o;
  wire n10326_o;
  wire n10327_o;
  wire n10328_o;
  wire n10332_o;
  wire n10333_o;
  wire [4:0] n10335_o;
  wire n10337_o;
  wire n10340_o;
  wire n10341_o;
  wire n10342_o;
  wire n10343_o;
  wire n10347_o;
  wire n10348_o;
  wire [4:0] n10350_o;
  wire n10352_o;
  wire n10355_o;
  wire n10356_o;
  wire n10357_o;
  wire n10358_o;
  wire n10362_o;
  wire n10363_o;
  wire [4:0] n10365_o;
  wire n10367_o;
  wire n10370_o;
  wire n10371_o;
  wire n10372_o;
  wire n10373_o;
  wire n10377_o;
  wire n10378_o;
  wire [4:0] n10380_o;
  wire n10382_o;
  wire n10385_o;
  wire n10386_o;
  wire n10387_o;
  wire n10388_o;
  wire n10392_o;
  wire n10393_o;
  wire [4:0] n10395_o;
  wire n10397_o;
  wire n10400_o;
  wire n10401_o;
  wire n10402_o;
  wire n10403_o;
  wire n10407_o;
  wire n10408_o;
  wire [4:0] n10410_o;
  wire n10412_o;
  wire n10415_o;
  wire n10416_o;
  wire n10417_o;
  wire n10418_o;
  wire n10422_o;
  wire n10423_o;
  wire [4:0] n10425_o;
  wire n10427_o;
  wire n10430_o;
  wire n10431_o;
  wire n10432_o;
  wire n10433_o;
  wire n10434_o;
  wire n10435_o;
  wire n10436_o;
  wire n10437_o;
  wire n10438_o;
  wire n10439_o;
  wire [4:0] n10440_o;
  wire n10442_o;
  wire n10445_o;
  wire n10446_o;
  wire [4:0] n10448_o;
  wire n10451_o;
  wire [31:0] n10452_o;
  wire [31:0] n10453_o;
  wire n10454_o;
  wire [15:0] n10455_o;
  wire [15:0] n10456_o;
  wire [31:0] n10457_o;
  wire [31:0] n10458_o;
  wire n10459_o;
  wire [23:0] n10460_o;
  wire [7:0] n10461_o;
  wire [31:0] n10462_o;
  wire [31:0] n10463_o;
  wire n10464_o;
  wire [35:0] n10466_o;
  wire [3:0] n10467_o;
  wire [3:0] n10468_o;
  wire [3:0] n10469_o;
  wire [31:0] n10470_o;
  wire [35:0] n10472_o;
  wire [35:0] n10473_o;
  wire [35:0] n10474_o;
  wire n10475_o;
  wire [37:0] n10477_o;
  wire [1:0] n10478_o;
  wire [1:0] n10479_o;
  wire [1:0] n10480_o;
  wire [35:0] n10481_o;
  wire [37:0] n10483_o;
  wire [37:0] n10484_o;
  wire [37:0] n10485_o;
  wire n10486_o;
  wire [38:0] n10488_o;
  wire [39:0] n10490_o;
  wire n10491_o;
  wire n10492_o;
  wire n10493_o;
  wire [38:0] n10494_o;
  wire [39:0] n10496_o;
  wire [39:0] n10497_o;
  wire [39:0] n10498_o;
  wire [39:0] n10499_o;
  wire [7:0] n10500_o;
  wire [7:0] n10501_o;
  wire [7:0] n10502_o;
  wire [31:0] n10503_o;
  wire n10504_o;
  wire n10505_o;
  wire [38:0] n10506_o;
  wire [39:0] n10507_o;
  wire [39:0] n10508_o;
  wire n10509_o;
  wire [1:0] n10510_o;
  wire [37:0] n10511_o;
  wire [39:0] n10512_o;
  wire [39:0] n10513_o;
  wire n10514_o;
  wire [3:0] n10515_o;
  wire [35:0] n10516_o;
  wire [39:0] n10517_o;
  wire [39:0] n10518_o;
  wire n10519_o;
  wire [7:0] n10520_o;
  wire [23:0] n10521_o;
  wire [31:0] n10522_o;
  wire [31:0] n10523_o;
  wire [31:0] n10524_o;
  wire n10525_o;
  wire [15:0] n10526_o;
  wire [15:0] n10527_o;
  wire [31:0] n10528_o;
  wire [31:0] n10529_o;
  wire [7:0] n10530_o;
  wire [31:0] n10531_o;
  wire [7:0] n10532_o;
  wire [39:0] n10533_o;
  localparam [39:0] n10534_o = 40'b0000000000000000000000000000000000000000;
  wire [39:0] n10536_o;
  localparam [39:0] n10538_o = 40'b1111111111111111111111111111111111111111;
  wire [39:0] n10540_o;
  wire [39:0] n10541_o;
  wire [39:0] n10542_o;
  wire n10543_o;
  wire n10544_o;
  wire n10545_o;
  wire n10546_o;
  wire n10547_o;
  wire n10548_o;
  wire n10549_o;
  wire n10550_o;
  wire n10551_o;
  wire n10552_o;
  wire n10560_o;
  wire n10561_o;
  wire n10562_o;
  wire n10563_o;
  wire n10564_o;
  wire n10565_o;
  wire n10566_o;
  wire n10567_o;
  wire n10568_o;
  wire n10569_o;
  wire n10577_o;
  wire n10578_o;
  wire n10579_o;
  wire n10580_o;
  wire n10581_o;
  wire n10582_o;
  wire n10583_o;
  wire n10584_o;
  wire n10585_o;
  wire n10586_o;
  wire n10594_o;
  wire n10595_o;
  wire n10596_o;
  wire n10597_o;
  wire n10598_o;
  wire n10599_o;
  wire n10600_o;
  wire n10601_o;
  wire n10602_o;
  wire n10603_o;
  wire n10611_o;
  wire n10612_o;
  wire n10613_o;
  wire n10614_o;
  wire n10615_o;
  wire n10616_o;
  wire n10617_o;
  wire n10618_o;
  wire n10619_o;
  wire n10620_o;
  wire n10628_o;
  wire n10629_o;
  wire n10630_o;
  wire n10631_o;
  wire n10632_o;
  wire n10633_o;
  wire n10634_o;
  wire n10635_o;
  wire n10636_o;
  wire n10637_o;
  wire n10645_o;
  wire n10646_o;
  wire n10647_o;
  wire n10648_o;
  wire n10649_o;
  wire n10650_o;
  wire n10651_o;
  wire n10652_o;
  wire n10653_o;
  wire n10654_o;
  wire n10662_o;
  wire n10663_o;
  wire n10664_o;
  wire n10665_o;
  wire n10666_o;
  wire n10667_o;
  wire n10668_o;
  wire n10669_o;
  wire n10670_o;
  wire n10671_o;
  wire n10679_o;
  wire n10680_o;
  wire n10681_o;
  wire n10682_o;
  wire n10683_o;
  wire n10684_o;
  wire n10685_o;
  wire n10686_o;
  wire n10687_o;
  wire n10688_o;
  wire n10696_o;
  wire n10697_o;
  wire n10698_o;
  wire n10699_o;
  wire n10700_o;
  wire n10701_o;
  wire n10702_o;
  wire n10703_o;
  wire n10704_o;
  wire n10705_o;
  wire n10713_o;
  wire n10714_o;
  wire n10715_o;
  wire n10716_o;
  wire n10717_o;
  wire n10718_o;
  wire n10719_o;
  wire n10720_o;
  wire n10721_o;
  wire n10722_o;
  wire n10730_o;
  wire n10731_o;
  wire n10732_o;
  wire n10733_o;
  wire n10734_o;
  wire n10735_o;
  wire n10736_o;
  wire n10737_o;
  wire n10738_o;
  wire n10739_o;
  wire n10747_o;
  wire n10748_o;
  wire n10749_o;
  wire n10750_o;
  wire n10751_o;
  wire n10752_o;
  wire n10753_o;
  wire n10754_o;
  wire n10755_o;
  wire n10756_o;
  wire n10764_o;
  wire n10765_o;
  wire n10766_o;
  wire n10767_o;
  wire n10768_o;
  wire n10769_o;
  wire n10770_o;
  wire n10771_o;
  wire n10772_o;
  wire n10773_o;
  wire n10781_o;
  wire n10782_o;
  wire n10783_o;
  wire n10784_o;
  wire n10785_o;
  wire n10786_o;
  wire n10787_o;
  wire n10788_o;
  wire n10789_o;
  wire n10790_o;
  wire n10798_o;
  wire n10799_o;
  wire n10800_o;
  wire n10801_o;
  wire n10802_o;
  wire n10803_o;
  wire n10804_o;
  wire n10805_o;
  wire n10806_o;
  wire n10807_o;
  wire n10815_o;
  wire n10816_o;
  wire n10817_o;
  wire n10818_o;
  wire n10819_o;
  wire n10820_o;
  wire n10821_o;
  wire n10822_o;
  wire n10823_o;
  wire n10824_o;
  wire n10832_o;
  wire n10833_o;
  wire n10834_o;
  wire n10835_o;
  wire n10836_o;
  wire n10837_o;
  wire n10838_o;
  wire n10839_o;
  wire n10840_o;
  wire n10841_o;
  wire n10849_o;
  wire n10850_o;
  wire n10851_o;
  wire n10852_o;
  wire n10853_o;
  wire n10854_o;
  wire n10855_o;
  wire n10856_o;
  wire n10857_o;
  wire n10858_o;
  wire n10866_o;
  wire n10867_o;
  wire n10868_o;
  wire n10869_o;
  wire n10870_o;
  wire n10871_o;
  wire n10872_o;
  wire n10873_o;
  wire n10874_o;
  wire n10875_o;
  wire n10883_o;
  wire n10884_o;
  wire n10885_o;
  wire n10886_o;
  wire n10887_o;
  wire n10888_o;
  wire n10889_o;
  wire n10890_o;
  wire n10891_o;
  wire n10892_o;
  wire n10900_o;
  wire n10901_o;
  wire n10902_o;
  wire n10903_o;
  wire n10904_o;
  wire n10905_o;
  wire n10906_o;
  wire n10907_o;
  wire n10908_o;
  wire n10909_o;
  wire n10917_o;
  wire n10918_o;
  wire n10919_o;
  wire n10920_o;
  wire n10921_o;
  wire n10922_o;
  wire n10923_o;
  wire n10924_o;
  wire n10925_o;
  wire n10926_o;
  wire n10934_o;
  wire n10935_o;
  wire n10936_o;
  wire n10937_o;
  wire n10938_o;
  wire n10939_o;
  wire n10940_o;
  wire n10941_o;
  wire n10942_o;
  wire n10943_o;
  wire n10951_o;
  wire n10952_o;
  wire n10953_o;
  wire n10954_o;
  wire n10955_o;
  wire n10956_o;
  wire n10957_o;
  wire n10958_o;
  wire n10959_o;
  wire n10960_o;
  wire n10968_o;
  wire n10969_o;
  wire n10970_o;
  wire n10971_o;
  wire n10972_o;
  wire n10973_o;
  wire n10974_o;
  wire n10975_o;
  wire n10976_o;
  wire n10977_o;
  wire n10985_o;
  wire n10986_o;
  wire n10987_o;
  wire n10988_o;
  wire n10989_o;
  wire n10990_o;
  wire n10991_o;
  wire n10992_o;
  wire n10993_o;
  wire n10994_o;
  wire n11002_o;
  wire n11003_o;
  wire n11004_o;
  wire n11005_o;
  wire n11006_o;
  wire n11007_o;
  wire n11008_o;
  wire n11009_o;
  wire n11010_o;
  wire n11011_o;
  wire n11019_o;
  wire n11020_o;
  wire n11021_o;
  wire n11022_o;
  wire n11023_o;
  wire n11024_o;
  wire n11025_o;
  wire n11026_o;
  wire n11027_o;
  wire n11028_o;
  wire n11036_o;
  wire n11037_o;
  wire n11038_o;
  wire n11039_o;
  wire n11040_o;
  wire n11041_o;
  wire n11042_o;
  wire n11043_o;
  wire n11044_o;
  wire n11045_o;
  wire n11053_o;
  wire n11054_o;
  wire n11055_o;
  wire n11056_o;
  wire n11057_o;
  wire n11058_o;
  wire n11059_o;
  wire n11060_o;
  wire n11061_o;
  wire n11062_o;
  wire n11070_o;
  wire n11071_o;
  wire n11072_o;
  wire n11073_o;
  wire n11074_o;
  wire n11075_o;
  wire n11076_o;
  wire n11077_o;
  wire n11078_o;
  wire n11079_o;
  wire n11087_o;
  wire n11088_o;
  wire n11089_o;
  wire n11090_o;
  wire n11091_o;
  wire n11092_o;
  wire n11093_o;
  wire n11094_o;
  wire n11095_o;
  wire n11096_o;
  wire n11104_o;
  wire n11105_o;
  wire n11106_o;
  wire n11107_o;
  wire n11108_o;
  wire n11109_o;
  wire n11110_o;
  wire n11111_o;
  wire n11112_o;
  wire n11113_o;
  wire n11121_o;
  wire n11122_o;
  wire n11123_o;
  wire n11124_o;
  wire n11125_o;
  wire n11126_o;
  wire n11127_o;
  wire n11128_o;
  wire n11129_o;
  wire n11130_o;
  wire n11138_o;
  wire n11139_o;
  wire n11140_o;
  wire n11141_o;
  wire n11142_o;
  wire n11143_o;
  wire n11144_o;
  wire n11145_o;
  wire n11146_o;
  wire n11147_o;
  wire n11155_o;
  wire n11156_o;
  wire n11157_o;
  wire n11158_o;
  wire n11159_o;
  wire n11160_o;
  wire n11161_o;
  wire n11162_o;
  wire n11163_o;
  wire n11164_o;
  wire n11172_o;
  wire n11173_o;
  wire n11174_o;
  wire n11175_o;
  wire n11176_o;
  wire n11177_o;
  wire n11178_o;
  wire n11179_o;
  wire n11180_o;
  wire n11181_o;
  wire n11189_o;
  wire n11190_o;
  wire n11191_o;
  wire n11192_o;
  wire n11193_o;
  wire n11194_o;
  wire n11195_o;
  wire n11196_o;
  wire n11197_o;
  wire n11198_o;
  wire n11199_o;
  wire n11200_o;
  wire n11201_o;
  wire n11202_o;
  wire n11203_o;
  wire n11204_o;
  wire n11205_o;
  wire n11206_o;
  wire n11207_o;
  wire n11208_o;
  wire [5:0] n11210_o;
  wire [5:0] n11211_o;
  wire [5:0] n11212_o;
  wire [3:0] n11213_o;
  wire n11215_o;
  wire [3:0] n11216_o;
  wire n11218_o;
  wire [3:0] n11219_o;
  wire n11221_o;
  wire [3:0] n11222_o;
  wire n11224_o;
  wire [3:0] n11226_o;
  wire n11228_o;
  wire [3:0] n11229_o;
  wire n11231_o;
  wire [3:0] n11233_o;
  wire n11235_o;
  wire [3:0] n11237_o;
  wire [3:0] n11238_o;
  wire [3:0] n11239_o;
  wire n11241_o;
  wire [3:0] n11242_o;
  wire [3:0] n11244_o;
  wire [1:0] n11245_o;
  wire n11246_o;
  wire n11247_o;
  wire n11248_o;
  wire n11250_o;
  wire [3:0] n11251_o;
  wire [3:0] n11252_o;
  wire [1:0] n11253_o;
  wire [1:0] n11255_o;
  wire [3:0] n11256_o;
  wire [3:0] n11259_o;
  wire [1:0] n11260_o;
  wire [2:0] n11261_o;
  wire [1:0] n11262_o;
  wire [1:0] n11263_o;
  wire n11264_o;
  wire n11266_o;
  wire [3:0] n11267_o;
  wire [3:0] n11269_o;
  wire [2:0] n11270_o;
  wire n11271_o;
  wire n11273_o;
  wire n11274_o;
  wire n11275_o;
  wire n11276_o;
  wire n11278_o;
  wire [3:0] n11279_o;
  wire [3:0] n11281_o;
  wire [2:0] n11282_o;
  wire n11283_o;
  wire n11284_o;
  wire [1:0] n11285_o;
  wire [1:0] n11287_o;
  wire [3:0] n11288_o;
  wire [3:0] n11289_o;
  wire [2:0] n11290_o;
  wire [2:0] n11292_o;
  localparam [4:0] n11293_o = 5'b11111;
  wire [1:0] n11295_o;
  wire n11297_o;
  wire n11299_o;
  wire n11300_o;
  wire n11302_o;
  wire n11303_o;
  wire n11306_o;
  wire n11307_o;
  wire n11308_o;
  wire n11310_o;
  wire n11311_o;
  wire n11312_o;
  wire n11314_o;
  wire n11315_o;
  wire [1:0] n11316_o;
  wire n11317_o;
  wire n11318_o;
  wire n11319_o;
  wire n11320_o;
  wire n11321_o;
  wire n11324_o;
  wire [1:0] n11329_o;
  wire n11330_o;
  wire n11332_o;
  wire n11333_o;
  wire n11335_o;
  wire n11337_o;
  wire n11338_o;
  wire n11339_o;
  wire n11341_o;
  wire [2:0] n11342_o;
  reg n11343_o;
  wire n11361_o;
  wire n11362_o;
  wire n11364_o;
  wire n11365_o;
  wire n11367_o;
  wire n11368_o;
  wire n11371_o;
  wire n11372_o;
  wire n11392_o;
  wire n11393_o;
  wire n11396_o;
  wire n11397_o;
  wire [31:0] n11398_o;
  wire n11403_o;
  wire [1:0] n11404_o;
  wire n11406_o;
  wire n11408_o;
  wire n11410_o;
  wire n11411_o;
  wire n11413_o;
  wire [2:0] n11414_o;
  reg [5:0] n11419_o;
  wire [1:0] n11420_o;
  wire n11422_o;
  wire n11424_o;
  wire n11426_o;
  wire n11427_o;
  wire n11429_o;
  wire [2:0] n11430_o;
  reg [5:0] n11435_o;
  wire [5:0] n11436_o;
  wire [1:0] n11438_o;
  wire n11440_o;
  wire n11441_o;
  wire n11442_o;
  wire n11443_o;
  wire n11444_o;
  wire [5:0] n11445_o;
  wire [2:0] n11446_o;
  wire [2:0] n11447_o;
  wire n11449_o;
  wire [2:0] n11452_o;
  wire [5:0] n11453_o;
  wire [5:0] n11454_o;
  wire [5:0] n11456_o;
  localparam [33:0] n11459_o = 34'b0000000000000000000000000000000000;
  wire n11463_o;
  wire [5:0] n11464_o;
  wire [5:0] n11466_o;
  wire [30:0] n11468_o;
  wire [31:0] n11470_o;
  wire [30:0] n11471_o;
  wire [31:0] n11473_o;
  wire [31:0] n11474_o;
  wire [32:0] n11475_o;
  wire [1:0] n11476_o;
  wire n11479_o;
  wire n11482_o;
  wire n11484_o;
  wire n11485_o;
  wire [1:0] n11486_o;
  wire n11487_o;
  reg n11488_o;
  wire n11489_o;
  reg n11490_o;
  wire [7:0] n11492_o;
  wire [15:0] n11493_o;
  wire [6:0] n11494_o;
  wire [31:0] n11495_o;
  wire [32:0] n11497_o;
  wire [32:0] n11498_o;
  wire n11500_o;
  wire n11501_o;
  wire n11502_o;
  wire n11503_o;
  wire n11504_o;
  wire n11506_o;
  wire n11508_o;
  wire n11509_o;
  wire n11510_o;
  wire [1:0] n11511_o;
  wire n11512_o;
  wire n11514_o;
  wire n11515_o;
  wire n11517_o;
  wire n11519_o;
  wire n11520_o;
  wire n11521_o;
  wire n11523_o;
  wire [2:0] n11524_o;
  reg n11525_o;
  wire n11526_o;
  wire n11528_o;
  wire n11529_o;
  wire [1:0] n11530_o;
  wire [7:0] n11531_o;
  wire [7:0] n11532_o;
  wire [7:0] n11533_o;
  wire n11534_o;
  wire n11536_o;
  wire [15:0] n11537_o;
  wire [15:0] n11538_o;
  wire [15:0] n11539_o;
  wire n11540_o;
  wire n11542_o;
  wire n11544_o;
  wire n11545_o;
  wire [31:0] n11546_o;
  wire [31:0] n11547_o;
  wire [31:0] n11548_o;
  wire n11549_o;
  wire n11551_o;
  wire [2:0] n11552_o;
  wire [7:0] n11553_o;
  wire [7:0] n11554_o;
  reg [7:0] n11556_o;
  wire [7:0] n11557_o;
  wire [7:0] n11558_o;
  reg [7:0] n11560_o;
  wire [15:0] n11561_o;
  reg [15:0] n11563_o;
  reg n11564_o;
  wire n11565_o;
  wire n11566_o;
  wire n11567_o;
  wire n11569_o;
  wire [1:0] n11570_o;
  wire [7:0] n11571_o;
  wire [7:0] n11572_o;
  wire [7:0] n11573_o;
  wire n11574_o;
  wire n11575_o;
  wire n11576_o;
  wire n11578_o;
  wire [15:0] n11579_o;
  wire [15:0] n11580_o;
  wire [15:0] n11581_o;
  wire n11582_o;
  wire n11583_o;
  wire n11584_o;
  wire n11586_o;
  wire n11588_o;
  wire n11589_o;
  wire [31:0] n11590_o;
  wire [31:0] n11591_o;
  wire [31:0] n11592_o;
  wire n11593_o;
  wire n11594_o;
  wire n11595_o;
  wire n11597_o;
  wire [2:0] n11598_o;
  wire [7:0] n11599_o;
  wire [7:0] n11600_o;
  reg [7:0] n11602_o;
  wire [7:0] n11603_o;
  wire [7:0] n11604_o;
  reg [7:0] n11606_o;
  wire [15:0] n11607_o;
  reg [15:0] n11609_o;
  reg n11610_o;
  wire n11611_o;
  wire n11612_o;
  wire [31:0] n11613_o;
  wire [31:0] n11614_o;
  wire [31:0] n11615_o;
  wire [31:0] n11616_o;
  wire [31:0] n11617_o;
  wire n11618_o;
  wire [31:0] n11619_o;
  wire [31:0] n11620_o;
  wire n11622_o;
  wire n11623_o;
  wire n11625_o;
  wire n11627_o;
  wire n11628_o;
  wire n11630_o;
  wire n11631_o;
  wire n11633_o;
  wire n11634_o;
  wire n11635_o;
  wire n11637_o;
  wire n11639_o;
  wire [5:0] n11641_o;
  wire n11643_o;
  wire [5:0] n11645_o;
  wire n11647_o;
  wire [5:0] n11649_o;
  wire n11651_o;
  wire [5:0] n11653_o;
  wire n11655_o;
  wire [5:0] n11657_o;
  wire n11659_o;
  wire [5:0] n11661_o;
  wire [5:0] n11662_o;
  wire [5:0] n11663_o;
  wire [5:0] n11664_o;
  wire [5:0] n11665_o;
  wire [5:0] n11666_o;
  wire [5:0] n11667_o;
  wire [5:0] n11669_o;
  wire n11671_o;
  wire n11673_o;
  wire [5:0] n11675_o;
  wire n11677_o;
  wire [5:0] n11679_o;
  wire n11681_o;
  wire [5:0] n11683_o;
  wire [5:0] n11684_o;
  wire [5:0] n11685_o;
  wire [5:0] n11686_o;
  wire n11688_o;
  wire n11690_o;
  wire [5:0] n11692_o;
  wire [5:0] n11693_o;
  wire n11695_o;
  wire [2:0] n11696_o;
  wire [5:0] n11698_o;
  wire n11700_o;
  wire [3:0] n11701_o;
  wire [5:0] n11703_o;
  wire n11705_o;
  wire [4:0] n11706_o;
  wire [5:0] n11708_o;
  wire n11710_o;
  wire [5:0] n11711_o;
  reg [5:0] n11713_o;
  wire n11714_o;
  wire n11715_o;
  wire [5:0] n11716_o;
  wire [5:0] n11717_o;
  wire n11718_o;
  wire n11719_o;
  wire n11720_o;
  wire n11721_o;
  wire [5:0] n11723_o;
  wire [5:0] n11724_o;
  wire n11725_o;
  wire n11726_o;
  wire n11727_o;
  wire [5:0] n11729_o;
  wire [5:0] n11730_o;
  wire [5:0] n11731_o;
  wire n11732_o;
  wire n11733_o;
  wire n11734_o;
  wire [5:0] n11736_o;
  wire [5:0] n11738_o;
  wire n11740_o;
  wire [5:0] n11741_o;
  wire n11742_o;
  wire [5:0] n11743_o;
  wire n11744_o;
  wire [31:0] n11745_o;
  wire [31:0] n11746_o;
  wire [31:0] n11747_o;
  localparam [32:0] n11748_o = 33'b000000000000000000000000000000000;
  wire n11749_o;
  wire n11751_o;
  wire n11752_o;
  wire n11753_o;
  wire n11754_o;
  wire n11755_o;
  wire [31:0] n11756_o;
  wire [31:0] n11757_o;
  wire n11758_o;
  wire n11760_o;
  wire n11762_o;
  wire [32:0] n11764_o;
  wire [1:0] n11765_o;
  wire n11766_o;
  localparam [23:0] n11767_o = 24'b000000000000000000000000;
  localparam [23:0] n11768_o = 24'b000000000000000000000000;
  wire n11770_o;
  wire n11771_o;
  wire n11772_o;
  wire n11773_o;
  wire [22:0] n11774_o;
  wire n11776_o;
  wire n11777_o;
  localparam [15:0] n11778_o = 16'b0000000000000000;
  wire n11781_o;
  wire n11782_o;
  wire n11783_o;
  wire n11784_o;
  wire [14:0] n11785_o;
  wire n11787_o;
  wire n11789_o;
  wire n11790_o;
  wire n11791_o;
  wire n11793_o;
  wire n11794_o;
  wire n11795_o;
  wire n11796_o;
  wire n11798_o;
  wire [2:0] n11799_o;
  wire n11800_o;
  reg n11801_o;
  wire [6:0] n11802_o;
  wire [6:0] n11803_o;
  reg [6:0] n11804_o;
  wire n11805_o;
  wire n11806_o;
  reg n11807_o;
  wire [14:0] n11808_o;
  wire [14:0] n11809_o;
  reg [14:0] n11810_o;
  wire n11811_o;
  reg n11812_o;
  wire [7:0] n11814_o;
  reg n11818_o;
  wire [7:0] n11819_o;
  wire [7:0] n11820_o;
  wire [7:0] n11821_o;
  wire [7:0] n11822_o;
  reg [7:0] n11823_o;
  wire [15:0] n11824_o;
  wire [15:0] n11825_o;
  wire [15:0] n11826_o;
  wire [15:0] n11827_o;
  reg [15:0] n11828_o;
  wire [7:0] n11832_o;
  wire [7:0] n11833_o;
  wire [7:0] n11834_o;
  wire [65:0] n11836_o;
  wire [30:0] n11837_o;
  wire [31:0] n11838_o;
  wire [65:0] n11839_o;
  wire n11843_o;
  wire [7:0] n11844_o;
  wire [7:0] n11845_o;
  wire n11846_o;
  wire [7:0] n11847_o;
  wire [7:0] n11848_o;
  wire n11849_o;
  wire [7:0] n11850_o;
  wire [7:0] n11851_o;
  wire [7:0] n11852_o;
  wire [7:0] n11853_o;
  wire [7:0] n11854_o;
  wire [7:0] n11855_o;
  wire n11856_o;
  wire n11857_o;
  wire n11858_o;
  wire n11859_o;
  wire [7:0] n11860_o;
  wire n11862_o;
  wire [7:0] n11864_o;
  wire n11866_o;
  wire [15:0] n11868_o;
  wire n11870_o;
  wire n11873_o;
  wire [1:0] n11874_o;
  wire [1:0] n11876_o;
  wire [2:0] n11877_o;
  wire [2:0] n11879_o;
  wire [2:0] n11881_o;
  wire n11884_o;
  wire n11885_o;
  wire n11886_o;
  wire [1:0] n11887_o;
  wire n11888_o;
  wire [2:0] n11889_o;
  wire n11890_o;
  wire [3:0] n11891_o;
  wire n11892_o;
  wire n11893_o;
  wire n11894_o;
  wire [1:0] n11895_o;
  wire [1:0] n11896_o;
  wire [1:0] n11897_o;
  wire [1:0] n11898_o;
  wire n11900_o;
  wire n11901_o;
  wire n11902_o;
  wire n11903_o;
  wire n11904_o;
  wire [1:0] n11905_o;
  wire n11906_o;
  wire [2:0] n11907_o;
  wire n11908_o;
  wire [3:0] n11909_o;
  wire n11910_o;
  wire n11911_o;
  wire [1:0] n11912_o;
  wire n11913_o;
  wire [2:0] n11914_o;
  wire n11915_o;
  wire [3:0] n11916_o;
  wire [3:0] n11917_o;
  wire [3:0] n11918_o;
  wire [3:0] n11919_o;
  wire n11921_o;
  wire n11922_o;
  wire n11925_o;
  wire n11928_o;
  wire n11929_o;
  wire n11930_o;
  wire n11931_o;
  wire n11932_o;
  wire n11933_o;
  wire n11935_o;
  wire n11936_o;
  wire n11938_o;
  wire n11939_o;
  wire n11940_o;
  wire n11941_o;
  wire n11942_o;
  wire [1:0] n11944_o;
  wire [3:0] n11946_o;
  wire [3:0] n11948_o;
  wire [3:0] n11949_o;
  wire [3:0] n11950_o;
  wire [3:0] n11951_o;
  wire [3:0] n11952_o;
  wire [3:0] n11953_o;
  wire [3:0] n11954_o;
  wire n11955_o;
  wire n11956_o;
  wire [3:0] n11957_o;
  wire n11958_o;
  wire n11959_o;
  wire n11960_o;
  wire n11962_o;
  wire n11963_o;
  wire n11964_o;
  wire n11965_o;
  wire n11966_o;
  wire n11967_o;
  wire n11968_o;
  wire n11969_o;
  wire n11970_o;
  wire n11971_o;
  wire n11972_o;
  wire n11973_o;
  wire n11974_o;
  wire n11975_o;
  wire n11976_o;
  wire n11977_o;
  wire n11978_o;
  wire n11979_o;
  wire n11981_o;
  wire n11983_o;
  wire n11985_o;
  wire n11986_o;
  wire n11987_o;
  wire [1:0] n11988_o;
  wire [3:0] n11990_o;
  wire n11991_o;
  wire n11992_o;
  wire [1:0] n11993_o;
  wire [3:0] n11995_o;
  wire [3:0] n11996_o;
  wire [3:0] n11997_o;
  wire n11998_o;
  wire n12000_o;
  wire n12001_o;
  wire n12002_o;
  wire n12003_o;
  wire n12004_o;
  wire n12007_o;
  wire n12009_o;
  wire n12010_o;
  wire n12011_o;
  wire n12013_o;
  wire n12014_o;
  wire n12015_o;
  wire n12016_o;
  wire n12017_o;
  wire n12018_o;
  wire n12019_o;
  wire n12020_o;
  wire n12021_o;
  wire n12022_o;
  wire n12023_o;
  wire n12024_o;
  wire n12025_o;
  wire n12026_o;
  wire n12028_o;
  wire n12029_o;
  wire n12032_o;
  wire n12033_o;
  wire n12034_o;
  wire n12035_o;
  wire n12036_o;
  wire [1:0] n12037_o;
  wire n12039_o;
  wire n12040_o;
  wire n12041_o;
  wire n12042_o;
  wire n12043_o;
  wire n12046_o;
  wire n12047_o;
  wire [1:0] n12048_o;
  wire n12049_o;
  wire n12050_o;
  wire n12051_o;
  wire n12052_o;
  wire n12053_o;
  wire n12054_o;
  wire n12055_o;
  wire n12056_o;
  wire n12057_o;
  wire n12058_o;
  wire n12059_o;
  wire n12060_o;
  wire n12061_o;
  wire n12062_o;
  wire n12063_o;
  wire n12064_o;
  wire n12065_o;
  wire n12066_o;
  wire n12067_o;
  wire n12068_o;
  wire n12069_o;
  wire n12070_o;
  wire n12072_o;
  wire n12073_o;
  wire n12074_o;
  wire n12075_o;
  wire n12076_o;
  wire n12077_o;
  wire n12079_o;
  wire n12080_o;
  wire n12081_o;
  wire n12082_o;
  wire [15:0] n12083_o;
  wire n12085_o;
  wire n12087_o;
  wire [15:0] n12088_o;
  wire n12090_o;
  wire n12091_o;
  wire n12092_o;
  wire n12095_o;
  wire [3:0] n12098_o;
  wire [3:0] n12099_o;
  wire [3:0] n12100_o;
  wire [3:0] n12101_o;
  wire [3:0] n12102_o;
  wire [3:0] n12103_o;
  wire [3:0] n12104_o;
  wire [3:0] n12105_o;
  wire [3:0] n12106_o;
  wire [1:0] n12107_o;
  wire [1:0] n12108_o;
  wire [1:0] n12109_o;
  wire [1:0] n12110_o;
  wire [1:0] n12111_o;
  wire [1:0] n12112_o;
  wire [1:0] n12113_o;
  wire n12114_o;
  wire n12115_o;
  wire n12116_o;
  wire n12117_o;
  wire n12118_o;
  wire n12119_o;
  wire n12120_o;
  wire n12121_o;
  wire n12122_o;
  wire [3:0] n12123_o;
  wire [3:0] n12124_o;
  wire [3:0] n12125_o;
  wire [3:0] n12126_o;
  wire [3:0] n12127_o;
  wire [3:0] n12128_o;
  wire [3:0] n12129_o;
  wire [3:0] n12130_o;
  wire [3:0] n12131_o;
  wire [3:0] n12132_o;
  wire [3:0] n12133_o;
  wire [3:0] n12134_o;
  wire [3:0] n12135_o;
  wire [4:0] n12136_o;
  wire [4:0] n12137_o;
  wire [4:0] n12138_o;
  wire [4:0] n12139_o;
  wire [4:0] n12140_o;
  wire [4:0] n12141_o;
  wire [4:0] n12142_o;
  wire [3:0] n12143_o;
  wire [3:0] n12144_o;
  wire [3:0] n12145_o;
  wire n12146_o;
  wire n12147_o;
  wire n12148_o;
  wire n12149_o;
  wire n12150_o;
  wire n12151_o;
  wire n12152_o;
  wire [3:0] n12153_o;
  wire [4:0] n12154_o;
  wire [4:0] n12155_o;
  wire [4:0] n12156_o;
  wire [2:0] n12157_o;
  wire [2:0] n12158_o;
  wire [2:0] n12159_o;
  wire [2:0] n12160_o;
  wire [2:0] n12161_o;
  wire [2:0] n12162_o;
  wire [2:0] n12163_o;
  wire [3:0] n12169_o;
  wire [7:0] n12170_o;
  wire [3:0] n12172_o;
  wire n12173_o;
  localparam [7:0] n12174_o = 8'b00000000;
  wire [3:0] n12176_o;
  wire n12177_o;
  wire [4:0] n12179_o;
  wire [4:0] n12180_o;
  wire [4:0] n12181_o;
  wire [4:0] n12182_o;
  wire [4:0] n12183_o;
  wire [7:0] n12184_o;
  wire n12191_o;
  wire n12192_o;
  wire n12193_o;
  wire [31:0] n12196_o;
  wire n12197_o;
  wire n12198_o;
  wire [31:0] n12201_o;
  wire [15:0] n12202_o;
  wire [15:0] n12203_o;
  wire n12204_o;
  wire n12205_o;
  wire [15:0] n12208_o;
  wire n12209_o;
  wire n12210_o;
  wire [15:0] n12213_o;
  wire [31:0] n12214_o;
  wire [31:0] n12215_o;
  wire [31:0] n12216_o;
  wire [31:0] n12217_o;
  wire [15:0] n12218_o;
  wire [47:0] n12219_o;
  wire [15:0] n12220_o;
  wire [63:0] n12221_o;
  wire [15:0] n12222_o;
  wire [47:0] n12223_o;
  wire [15:0] n12224_o;
  wire [63:0] n12225_o;
  wire [127:0] n12226_o;
  wire [127:0] n12227_o;
  wire [127:0] n12228_o;
  wire [31:0] n12229_o;
  wire n12231_o;
  wire n12232_o;
  wire n12233_o;
  wire n12234_o;
  wire n12235_o;
  wire n12236_o;
  wire [31:0] n12237_o;
  wire n12239_o;
  wire n12240_o;
  wire n12241_o;
  wire n12242_o;
  wire n12243_o;
  wire n12246_o;
  wire [31:0] n12251_o;
  wire n12259_o;
  wire n12260_o;
  wire n12261_o;
  wire n12262_o;
  wire n12263_o;
  wire n12264_o;
  wire n12265_o;
  wire n12266_o;
  wire n12268_o;
  wire n12269_o;
  wire n12270_o;
  wire n12271_o;
  wire n12272_o;
  wire n12273_o;
  wire n12274_o;
  wire n12275_o;
  wire n12276_o;
  wire n12277_o;
  wire n12278_o;
  wire n12279_o;
  wire n12280_o;
  wire n12281_o;
  wire n12282_o;
  wire n12283_o;
  wire n12284_o;
  wire n12285_o;
  wire n12286_o;
  wire n12287_o;
  wire n12288_o;
  wire n12289_o;
  wire n12290_o;
  wire n12291_o;
  wire n12292_o;
  wire n12293_o;
  wire n12294_o;
  wire n12295_o;
  wire n12296_o;
  wire n12297_o;
  wire n12298_o;
  wire n12299_o;
  wire n12300_o;
  wire n12301_o;
  wire n12302_o;
  wire n12303_o;
  wire n12304_o;
  wire n12305_o;
  wire n12306_o;
  wire n12307_o;
  wire n12308_o;
  wire n12309_o;
  wire n12310_o;
  wire n12311_o;
  wire n12312_o;
  wire n12313_o;
  wire n12314_o;
  wire n12315_o;
  wire n12316_o;
  wire n12317_o;
  wire n12318_o;
  wire n12319_o;
  wire n12320_o;
  wire n12321_o;
  wire n12322_o;
  wire n12323_o;
  wire n12324_o;
  wire n12325_o;
  wire n12326_o;
  wire n12327_o;
  wire n12328_o;
  wire n12329_o;
  wire n12330_o;
  wire n12331_o;
  wire [3:0] n12332_o;
  wire [3:0] n12333_o;
  wire [3:0] n12334_o;
  wire [3:0] n12335_o;
  wire [3:0] n12336_o;
  wire [3:0] n12337_o;
  wire [3:0] n12338_o;
  wire [3:0] n12339_o;
  wire [15:0] n12340_o;
  wire [15:0] n12341_o;
  wire [31:0] n12342_o;
  wire n12343_o;
  wire n12345_o;
  wire n12346_o;
  wire n12347_o;
  wire n12348_o;
  wire n12349_o;
  wire [31:0] n12350_o;
  wire n12351_o;
  wire n12352_o;
  wire [63:0] n12353_o;
  wire [15:0] n12354_o;
  wire [15:0] n12355_o;
  wire [31:0] n12356_o;
  wire [31:0] n12357_o;
  wire [15:0] n12358_o;
  wire [15:0] n12359_o;
  wire [15:0] n12360_o;
  wire n12362_o;
  wire n12363_o;
  wire n12364_o;
  wire [15:0] n12365_o;
  wire [15:0] n12367_o;
  wire n12368_o;
  wire n12369_o;
  wire [32:0] n12370_o;
  wire [32:0] n12372_o;
  wire [32:0] n12373_o;
  wire [32:0] n12374_o;
  wire [16:0] n12376_o;
  wire [15:0] n12377_o;
  wire [32:0] n12378_o;
  wire [32:0] n12379_o;
  wire [32:0] n12380_o;
  wire n12381_o;
  wire [31:0] n12382_o;
  wire [31:0] n12383_o;
  wire [31:0] n12384_o;
  wire [30:0] n12385_o;
  wire n12386_o;
  wire [31:0] n12387_o;
  wire [31:0] n12388_o;
  wire [31:0] n12390_o;
  wire [31:0] n12391_o;
  wire [31:0] n12392_o;
  wire n12393_o;
  wire n12394_o;
  wire n12395_o;
  wire n12396_o;
  wire n12397_o;
  wire n12398_o;
  wire n12399_o;
  wire n12400_o;
  wire n12401_o;
  wire n12402_o;
  wire n12403_o;
  wire n12404_o;
  wire n12406_o;
  wire n12409_o;
  wire n12415_o;
  wire n12418_o;
  wire n12419_o;
  wire n12420_o;
  wire [63:0] n12422_o;
  wire [63:0] n12423_o;
  wire n12426_o;
  wire n12427_o;
  wire n12428_o;
  wire [63:0] n12429_o;
  wire n12431_o;
  wire n12434_o;
  wire n12435_o;
  wire n12436_o;
  wire n12437_o;
  wire [31:0] n12438_o;
  wire [32:0] n12440_o;
  wire [16:0] n12442_o;
  wire [15:0] n12443_o;
  wire [32:0] n12444_o;
  wire [32:0] n12445_o;
  wire n12448_o;
  wire n12449_o;
  wire [31:0] n12450_o;
  wire [31:0] n12452_o;
  wire [31:0] n12453_o;
  wire [31:0] n12454_o;
  wire [63:0] n12455_o;
  wire n12457_o;
  wire n12458_o;
  wire n12460_o;
  wire n12461_o;
  wire n12464_o;
  wire [31:0] n12474_o;
  wire [2:0] n12475_o;
  wire [3:0] n12476_o;
  reg [3:0] n12477_q;
  wire [8:0] n12478_o;
  wire [63:0] n12479_o;
  reg [63:0] n12480_q;
  wire n12481_o;
  reg n12482_q;
  reg n12483_q;
  wire n12485_o;
  reg n12486_q;
  wire n12487_o;
  reg n12488_q;
  wire [31:0] n12492_o;
  wire [31:0] n12493_o;
  reg [31:0] n12494_q;
  wire [63:0] n12496_o;
  wire [63:0] n12498_o;
  reg [63:0] n12499_q;
  wire [63:0] n12500_o;
  wire n12502_o;
  reg n12503_q;
  wire [32:0] n12504_o;
  reg [32:0] n12505_q;
  wire n12506_o;
  reg n12507_q;
  wire [63:0] n12508_o;
  wire n12509_o;
  reg n12510_q;
  wire n12511_o;
  reg n12512_q;
  wire [31:0] n12515_o;
  wire [39:0] n12517_o;
  wire [31:0] n12518_o;
  wire [39:0] n12520_o;
  wire [4:0] n12521_o;
  wire n12522_o;
  reg n12523_q;
  wire n12524_o;
  reg n12525_q;
  wire n12526_o;
  reg n12527_q;
  wire n12528_o;
  reg n12529_q;
  wire n12530_o;
  reg n12531_q;
  wire n12532_o;
  reg n12533_q;
  wire n12534_o;
  reg n12535_q;
  wire [32:0] n12537_o;
  wire [32:0] n12538_o;
  wire [32:0] n12539_o;
  wire [31:0] n12540_o;
  wire [7:0] n12541_o;
  reg [7:0] n12542_q;
  reg [7:0] n12543_q;
  wire n12544_o;
  wire n12545_o;
  wire n12546_o;
  wire n12547_o;
  wire n12548_o;
  wire n12549_o;
  wire n12550_o;
  wire n12551_o;
  wire n12552_o;
  wire n12553_o;
  wire n12554_o;
  wire n12555_o;
  wire n12556_o;
  wire n12557_o;
  wire n12558_o;
  wire n12559_o;
  wire n12560_o;
  wire n12561_o;
  wire n12562_o;
  wire n12563_o;
  wire n12564_o;
  wire n12565_o;
  wire n12566_o;
  wire n12567_o;
  wire n12568_o;
  wire n12569_o;
  wire n12570_o;
  wire n12571_o;
  wire n12572_o;
  wire n12573_o;
  wire n12574_o;
  wire n12575_o;
  wire [1:0] n12576_o;
  reg n12577_o;
  wire [1:0] n12578_o;
  reg n12579_o;
  wire [1:0] n12580_o;
  reg n12581_o;
  wire [1:0] n12582_o;
  reg n12583_o;
  wire [1:0] n12584_o;
  reg n12585_o;
  wire [1:0] n12586_o;
  reg n12587_o;
  wire [1:0] n12588_o;
  reg n12589_o;
  wire [1:0] n12590_o;
  reg n12591_o;
  wire [1:0] n12592_o;
  reg n12593_o;
  wire [1:0] n12594_o;
  reg n12595_o;
  wire n12596_o;
  wire n12597_o;
  wire n12598_o;
  wire n12599_o;
  wire n12600_o;
  wire n12601_o;
  wire n12602_o;
  wire n12603_o;
  wire n12604_o;
  wire n12605_o;
  wire n12606_o;
  wire n12607_o;
  wire n12608_o;
  wire n12609_o;
  wire n12610_o;
  wire n12611_o;
  wire n12612_o;
  wire n12613_o;
  wire n12614_o;
  wire n12615_o;
  wire n12616_o;
  wire n12617_o;
  wire n12618_o;
  wire n12619_o;
  wire n12620_o;
  wire n12621_o;
  wire n12622_o;
  wire n12623_o;
  wire n12624_o;
  wire n12625_o;
  wire n12626_o;
  wire n12627_o;
  wire n12628_o;
  wire n12629_o;
  wire n12630_o;
  wire n12631_o;
  wire n12632_o;
  wire n12633_o;
  wire n12634_o;
  wire n12635_o;
  wire n12636_o;
  wire n12637_o;
  wire n12638_o;
  wire n12639_o;
  wire n12640_o;
  wire n12641_o;
  wire n12642_o;
  wire n12643_o;
  wire n12644_o;
  wire n12645_o;
  wire n12646_o;
  wire n12647_o;
  wire n12648_o;
  wire n12649_o;
  wire n12650_o;
  wire n12651_o;
  wire n12652_o;
  wire n12653_o;
  wire n12654_o;
  wire n12655_o;
  wire n12656_o;
  wire n12657_o;
  wire n12658_o;
  wire n12659_o;
  wire n12660_o;
  wire n12661_o;
  wire n12662_o;
  wire n12663_o;
  wire n12664_o;
  wire n12665_o;
  wire n12666_o;
  wire n12667_o;
  wire n12668_o;
  wire n12669_o;
  wire n12670_o;
  wire n12671_o;
  wire n12672_o;
  wire n12673_o;
  wire n12674_o;
  wire n12675_o;
  wire n12676_o;
  wire n12677_o;
  wire n12678_o;
  wire n12679_o;
  wire n12680_o;
  wire n12681_o;
  wire n12682_o;
  wire n12683_o;
  wire n12684_o;
  wire n12685_o;
  wire n12686_o;
  wire n12687_o;
  wire n12688_o;
  wire n12689_o;
  wire n12690_o;
  wire n12691_o;
  wire n12692_o;
  wire n12693_o;
  wire n12694_o;
  wire n12695_o;
  wire n12696_o;
  wire n12697_o;
  wire n12698_o;
  wire n12699_o;
  wire n12700_o;
  wire n12701_o;
  wire n12702_o;
  wire n12703_o;
  wire n12704_o;
  wire n12705_o;
  wire n12706_o;
  wire n12707_o;
  wire n12708_o;
  wire n12709_o;
  wire n12710_o;
  wire n12711_o;
  wire n12712_o;
  wire n12713_o;
  wire n12714_o;
  wire n12715_o;
  wire n12716_o;
  wire n12717_o;
  wire n12718_o;
  wire n12719_o;
  wire n12720_o;
  wire n12721_o;
  wire n12722_o;
  wire n12723_o;
  wire n12724_o;
  wire n12725_o;
  wire n12726_o;
  wire n12727_o;
  wire n12728_o;
  wire n12729_o;
  wire n12730_o;
  wire n12731_o;
  wire [31:0] n12732_o;
  wire n12733_o;
  wire n12734_o;
  wire n12735_o;
  wire n12736_o;
  wire n12737_o;
  wire n12738_o;
  wire n12739_o;
  wire n12740_o;
  wire n12741_o;
  wire n12742_o;
  wire n12743_o;
  wire n12744_o;
  wire n12745_o;
  wire n12746_o;
  wire n12747_o;
  wire n12748_o;
  wire n12749_o;
  wire n12750_o;
  wire n12751_o;
  wire n12752_o;
  wire n12753_o;
  wire n12754_o;
  wire n12755_o;
  wire n12756_o;
  wire n12757_o;
  wire n12758_o;
  wire n12759_o;
  wire n12760_o;
  wire n12761_o;
  wire n12762_o;
  wire n12763_o;
  wire n12764_o;
  wire [1:0] n12765_o;
  reg n12766_o;
  wire [1:0] n12767_o;
  reg n12768_o;
  wire [1:0] n12769_o;
  reg n12770_o;
  wire [1:0] n12771_o;
  reg n12772_o;
  wire [1:0] n12773_o;
  reg n12774_o;
  wire [1:0] n12775_o;
  reg n12776_o;
  wire [1:0] n12777_o;
  reg n12778_o;
  wire [1:0] n12779_o;
  reg n12780_o;
  wire [1:0] n12781_o;
  reg n12782_o;
  wire [1:0] n12783_o;
  reg n12784_o;
  wire n12785_o;
  wire n12786_o;
  wire n12787_o;
  wire n12788_o;
  wire n12789_o;
  wire n12790_o;
  wire n12791_o;
  wire n12792_o;
  wire n12793_o;
  wire n12794_o;
  wire n12795_o;
  wire n12796_o;
  wire n12797_o;
  wire n12798_o;
  wire n12799_o;
  wire n12800_o;
  wire n12801_o;
  wire n12802_o;
  wire n12803_o;
  wire n12804_o;
  wire n12805_o;
  wire n12806_o;
  wire n12807_o;
  wire n12808_o;
  wire n12809_o;
  wire n12810_o;
  wire n12811_o;
  wire n12812_o;
  wire n12813_o;
  wire n12814_o;
  wire n12815_o;
  wire n12816_o;
  wire n12817_o;
  wire n12818_o;
  wire n12819_o;
  wire n12820_o;
  wire n12821_o;
  wire n12822_o;
  wire n12823_o;
  wire n12824_o;
  wire n12825_o;
  wire n12826_o;
  wire n12827_o;
  wire n12828_o;
  wire n12829_o;
  wire n12830_o;
  wire n12831_o;
  wire n12832_o;
  wire n12833_o;
  wire n12834_o;
  wire n12835_o;
  wire n12836_o;
  wire n12837_o;
  wire n12838_o;
  wire n12839_o;
  wire n12840_o;
  wire n12841_o;
  wire n12842_o;
  wire n12843_o;
  wire n12844_o;
  wire n12845_o;
  wire n12846_o;
  wire n12847_o;
  wire n12848_o;
  wire n12849_o;
  wire n12850_o;
  wire n12851_o;
  wire n12852_o;
  wire n12853_o;
  wire n12854_o;
  wire n12855_o;
  wire n12856_o;
  wire n12857_o;
  wire n12858_o;
  wire n12859_o;
  wire n12860_o;
  wire n12861_o;
  wire n12862_o;
  wire n12863_o;
  wire n12864_o;
  wire n12865_o;
  wire n12866_o;
  wire n12867_o;
  wire n12868_o;
  wire n12869_o;
  wire n12870_o;
  wire n12871_o;
  wire n12872_o;
  wire n12873_o;
  wire n12874_o;
  wire n12875_o;
  wire n12876_o;
  wire n12877_o;
  wire n12878_o;
  wire n12879_o;
  wire n12880_o;
  wire n12881_o;
  wire n12882_o;
  wire n12883_o;
  wire n12884_o;
  wire n12885_o;
  wire n12886_o;
  wire n12887_o;
  wire n12888_o;
  wire n12889_o;
  wire n12890_o;
  wire n12891_o;
  wire n12892_o;
  wire n12893_o;
  wire n12894_o;
  wire n12895_o;
  wire n12896_o;
  wire n12897_o;
  wire n12898_o;
  wire n12899_o;
  wire n12900_o;
  wire n12901_o;
  wire n12902_o;
  wire n12903_o;
  wire n12904_o;
  wire n12905_o;
  wire n12906_o;
  wire n12907_o;
  wire n12908_o;
  wire n12909_o;
  wire n12910_o;
  wire n12911_o;
  wire n12912_o;
  wire n12913_o;
  wire n12914_o;
  wire n12915_o;
  wire n12916_o;
  wire n12917_o;
  wire n12918_o;
  wire n12919_o;
  wire n12920_o;
  wire n12921_o;
  wire n12922_o;
  wire n12923_o;
  wire n12924_o;
  wire n12925_o;
  wire n12926_o;
  wire n12927_o;
  wire n12928_o;
  wire n12929_o;
  wire n12930_o;
  wire n12931_o;
  wire n12932_o;
  wire n12933_o;
  wire n12934_o;
  wire [33:0] n12935_o;
  assign bf_ext_out = n12542_q;
  assign set_v_flag = n12409_o;
  assign flags = n12543_q;
  assign c_out = n9786_o;
  assign addsub_q = n9764_o;
  assign aluout = n9546_o;
  /* ../TG68K.C/TG68K_ALU.vhd:86:16  */
  assign op1in = n12474_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:87:16  */
  assign addsub_a = n9652_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:88:16  */
  assign addsub_b = n9735_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:89:16  */
  assign notaddsub_b = n9747_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:90:16  */
  assign add_result = n9752_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:91:16  */
  assign addsub_ofl = n12475_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:92:16  */
  assign opaddsub = n9714_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:93:16  */
  assign c_in = n12476_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:94:16  */
  assign flag_z = n11881_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:95:16  */
  assign set_flags = n11919_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:1013:67  */
  assign ccrin = n11855_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:97:16  */
  assign last_flags1 = n12477_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:100:16  */
  assign bcd_pur = n9792_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:101:16  */
  assign bcd_kor = n12478_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:102:16  */
  assign halve_carry = n9797_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:103:16  */
  assign vflag_a = n9850_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:104:16  */
  assign bcd_a_carry = n9853_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:105:16  */
  assign bcd_a = n9847_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:106:16  */
  assign result_mulu = n12228_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:107:16  */
  assign result_div = n12480_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:108:16  */
  assign result_div_pre = n12392_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:109:16  */
  assign set_mv_flag = n12246_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:110:16  */
  assign v_flag = n12482_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:112:16  */
  assign rot_rot = n11343_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:115:16  */
  assign rot_x = n11396_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:116:16  */
  assign rot_c = n11397_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:117:16  */
  assign rot_out = n11398_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:118:16  */
  assign asl_vflag = n12483_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:120:16  */
  assign bit_number = n9894_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:121:16  */
  assign bits_out = n12732_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:122:16  */
  assign one_bit_in = n12597_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:123:16  */
  assign bchg = n12486_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:124:16  */
  assign bset = n12488_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:129:16  */
  assign mulu_reg = n12496_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:1153:86  */
  assign faktora = n12215_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:1153:157  */
  assign faktorb = n12217_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:134:16  */
  assign div_reg = n12499_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:135:16  */
  assign div_quot = n12500_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:137:16  */
  assign div_neg = n12503_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:138:16  */
  assign div_bit = n12381_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:139:16  */
  assign div_sub = n12380_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:140:16  */
  assign div_over = n12505_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:141:16  */
  assign nozero = n12507_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:142:16  */
  assign div_qsign = n12352_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:143:16  */
  assign dividend = n12508_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:144:16  */
  assign divs = n12266_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:145:16  */
  assign signedop = n12510_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:146:16  */
  assign op1_sign = n12512_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:1316:103  */
  assign op2outext = n12367_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:151:16  */
  assign datareg = n12515_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:153:16  */
  assign bf_datareg = n10453_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:154:16  */
  assign result = n12517_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:155:16  */
  assign result_tmp = n10542_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:156:16  */
  assign unshifted_bitmask = n12518_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:158:16  */
  assign inmux0 = n10508_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:159:16  */
  assign inmux1 = n10513_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:160:16  */
  assign inmux2 = n10518_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:161:16  */
  assign inmux3 = n10524_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:162:16  */
  assign shifted_bitmask = n10498_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:163:16  */
  assign bitmaskmux0 = n10485_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:164:16  */
  assign bitmaskmux1 = n10474_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:165:16  */
  assign bitmaskmux2 = n10463_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:166:16  */
  assign bitmaskmux3 = n10458_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:167:16  */
  assign bf_set2 = n10529_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:168:16  */
  assign shift = n12520_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:169:16  */
  assign bf_firstbit = n11212_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:170:16  */
  assign mux = n11289_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:171:16  */
  assign bitnr = n12521_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:172:16  */
  assign mask = datareg; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:173:16  */
  assign mask_not_zero = n11324_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:174:16  */
  assign bf_bset = n12523_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:175:16  */
  assign bf_nflag = n12786_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:176:16  */
  assign bf_bchg = n12525_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:177:16  */
  assign bf_ins = n12527_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:178:16  */
  assign bf_exts = n12529_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:179:16  */
  assign bf_fffo = n12531_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:180:16  */
  assign bf_d32 = n12533_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:181:16  */
  assign bf_s32 = n12535_q; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:187:16  */
  assign hot_msb = n12935_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:188:16  */
  assign vector = n12537_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:189:16  */
  assign result_bs = n11839_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:946:110  */
  assign bit_nr = n11743_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:191:16  */
  assign bit_msb = n11466_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:192:16  */
  assign bs_shift = n11456_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:887:39  */
  assign bs_shift_mod = n11713_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:194:16  */
  assign asl_over = n11498_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:195:16  */
  assign asl_over_xor = n12538_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:196:16  */
  assign asr_sign = n12539_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:197:16  */
  assign msb = n11818_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:198:16  */
  assign ring = n11436_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:199:16  */
  assign alu = n11620_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:200:16  */
  assign bsout = n12540_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:201:16  */
  assign bs_v = n11633_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:202:16  */
  assign bs_c = n11760_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:203:16  */
  assign bs_x = n11635_o; // (signal)
  /* ../TG68K.C/TG68K_ALU.vhd:215:35  */
  assign n9536_o = op1in[7];
  /* ../TG68K.C/TG68K_ALU.vhd:215:39  */
  assign n9537_o = n9536_o | exec_tas;
  assign n9538_o = op1in[31:8];
  assign n9539_o = op1in[6:0];
  /* ../TG68K.C/TG68K_ALU.vhd:216:24  */
  assign n9540_o = exec[76];
  /* ../TG68K.C/TG68K_ALU.vhd:217:41  */
  assign n9541_o = result[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:219:57  */
  assign n9542_o = {26'b0, bf_firstbit};  //  uext
  /* ../TG68K.C/TG68K_ALU.vhd:219:57  */
  assign n9543_o = bf_ffo_offset - n9542_o;
  /* ../TG68K.C/TG68K_ALU.vhd:218:25  */
  assign n9544_o = bf_fffo ? n9543_o : n9541_o;
  assign n9545_o = {n9538_o, n9537_o, n9539_o};
  /* ../TG68K.C/TG68K_ALU.vhd:216:17  */
  assign n9546_o = n9540_o ? n9544_o : n9545_o;
  /* ../TG68K.C/TG68K_ALU.vhd:224:24  */
  assign n9547_o = exec[12];
  /* ../TG68K.C/TG68K_ALU.vhd:224:45  */
  assign n9548_o = exec[13];
  /* ../TG68K.C/TG68K_ALU.vhd:224:38  */
  assign n9549_o = n9547_o | n9548_o;
  /* ../TG68K.C/TG68K_ALU.vhd:225:51  */
  assign n9550_o = bcd_a[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:226:27  */
  assign n9551_o = exec[20];
  /* ../TG68K.C/TG68K_ALU.vhd:226:41  */
  assign n9553_o = n9551_o & 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:234:40  */
  assign n9554_o = exec[67];
  /* ../TG68K.C/TG68K_ALU.vhd:235:61  */
  assign n9555_o = result_mulu[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:238:58  */
  assign n9556_o = mulu_reg[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:234:33  */
  assign n9557_o = n9554_o ? n9555_o : n9556_o;
  /* ../TG68K.C/TG68K_ALU.vhd:241:27  */
  assign n9558_o = exec[21];
  /* ../TG68K.C/TG68K_ALU.vhd:241:41  */
  assign n9560_o = n9558_o & 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:242:38  */
  assign n9561_o = exe_opcode[15];
  /* ../TG68K.C/TG68K_ALU.vhd:242:47  */
  assign n9563_o = n9561_o | 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:244:52  */
  assign n9564_o = result_div[47:32];
  /* ../TG68K.C/TG68K_ALU.vhd:244:77  */
  assign n9565_o = result_div[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:244:66  */
  assign n9566_o = {n9564_o, n9565_o};
  /* ../TG68K.C/TG68K_ALU.vhd:246:40  */
  assign n9567_o = exec[68];
  /* ../TG68K.C/TG68K_ALU.vhd:247:60  */
  assign n9568_o = result_div[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:249:60  */
  assign n9569_o = result_div[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:246:33  */
  assign n9570_o = n9567_o ? n9568_o : n9569_o;
  /* ../TG68K.C/TG68K_ALU.vhd:242:25  */
  assign n9571_o = n9563_o ? n9566_o : n9570_o;
  /* ../TG68K.C/TG68K_ALU.vhd:252:27  */
  assign n9572_o = exec[5];
  /* ../TG68K.C/TG68K_ALU.vhd:253:41  */
  assign n9573_o = op2out | op1out;
  /* ../TG68K.C/TG68K_ALU.vhd:254:27  */
  assign n9574_o = exec[6];
  /* ../TG68K.C/TG68K_ALU.vhd:255:41  */
  assign n9575_o = op2out & op1out;
  /* ../TG68K.C/TG68K_ALU.vhd:256:27  */
  assign n9576_o = exec[16];
  assign n9577_o = {exe_condition, exe_condition, exe_condition, exe_condition};
  assign n9578_o = {exe_condition, exe_condition, exe_condition, exe_condition};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3097:71  */
  assign n9579_o = {n9577_o, n9578_o};
  /* ../TG68K.C/TG68K_ALU.vhd:258:27  */
  assign n9580_o = exec[7];
  /* ../TG68K.C/TG68K_ALU.vhd:259:41  */
  assign n9581_o = op2out ^ op1out;
  /* ../TG68K.C/TG68K_ALU.vhd:261:27  */
  assign n9582_o = exec[85];
  /* ../TG68K.C/TG68K_ALU.vhd:264:27  */
  assign n9583_o = exec[9];
  /* ../TG68K.C/TG68K_ALU.vhd:266:27  */
  assign n9584_o = exec[81];
  /* ../TG68K.C/TG68K_ALU.vhd:268:27  */
  assign n9585_o = exec[15];
  /* ../TG68K.C/TG68K_ALU.vhd:269:40  */
  assign n9586_o = op1out[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:269:61  */
  assign n9587_o = op1out[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:269:53  */
  assign n9588_o = {n9586_o, n9587_o};
  /* ../TG68K.C/TG68K_ALU.vhd:270:27  */
  assign n9589_o = exec[14];
  /* ../TG68K.C/TG68K_ALU.vhd:272:27  */
  assign n9590_o = exec[75];
  /* ../TG68K.C/TG68K_ALU.vhd:274:27  */
  assign n9591_o = exec[2];
  /* ../TG68K.C/TG68K_ALU.vhd:276:38  */
  assign n9592_o = exe_opcode[9];
  /* ../TG68K.C/TG68K_ALU.vhd:276:25  */
  assign n9594_o = n9592_o ? 8'b00000000 : flagssr;
  /* ../TG68K.C/TG68K_ALU.vhd:281:27  */
  assign n9595_o = exec[77];
  /* ../TG68K.C/TG68K_ALU.vhd:282:54  */
  assign n9596_o = n9764_o[11:8];
  /* ../TG68K.C/TG68K_ALU.vhd:282:78  */
  assign n9597_o = n9764_o[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:282:68  */
  assign n9598_o = {n9596_o, n9597_o};
  assign n9599_o = n9764_o[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:281:17  */
  assign n9600_o = n9595_o ? n9598_o : n9599_o;
  assign n9601_o = {n9594_o, n12543_q};
  assign n9602_o = n9601_o[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:274:17  */
  assign n9603_o = n9591_o ? n9602_o : n9600_o;
  assign n9604_o = n9601_o[15:8];
  assign n9605_o = n9764_o[15:8];
  /* ../TG68K.C/TG68K_ALU.vhd:274:17  */
  assign n9606_o = n9591_o ? n9604_o : n9605_o;
  assign n9607_o = {n9606_o, n9603_o};
  assign n9608_o = bf_datareg[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:272:17  */
  assign n9609_o = n9590_o ? n9608_o : n9607_o;
  assign n9610_o = bf_datareg[31:16];
  assign n9611_o = n9764_o[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:272:17  */
  assign n9612_o = n9590_o ? n9610_o : n9611_o;
  assign n9613_o = {n9612_o, n9609_o};
  /* ../TG68K.C/TG68K_ALU.vhd:270:17  */
  assign n9614_o = n9589_o ? bits_out : n9613_o;
  /* ../TG68K.C/TG68K_ALU.vhd:268:17  */
  assign n9615_o = n9585_o ? n9588_o : n9614_o;
  /* ../TG68K.C/TG68K_ALU.vhd:266:17  */
  assign n9616_o = n9584_o ? bsout : n9615_o;
  /* ../TG68K.C/TG68K_ALU.vhd:264:17  */
  assign n9617_o = n9583_o ? rot_out : n9616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:261:17  */
  assign n9618_o = n9582_o ? op2out : n9617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:258:17  */
  assign n9619_o = n9580_o ? n9581_o : n9618_o;
  assign n9620_o = n9619_o[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:256:17  */
  assign n9621_o = n9576_o ? n9579_o : n9620_o;
  assign n9622_o = n9619_o[31:8];
  assign n9623_o = n9764_o[31:8];
  /* ../TG68K.C/TG68K_ALU.vhd:256:17  */
  assign n9624_o = n9576_o ? n9623_o : n9622_o;
  assign n9625_o = {n9624_o, n9621_o};
  /* ../TG68K.C/TG68K_ALU.vhd:254:17  */
  assign n9626_o = n9574_o ? n9575_o : n9625_o;
  /* ../TG68K.C/TG68K_ALU.vhd:252:17  */
  assign n9627_o = n9572_o ? n9573_o : n9626_o;
  /* ../TG68K.C/TG68K_ALU.vhd:241:17  */
  assign n9628_o = n9560_o ? n9571_o : n9627_o;
  /* ../TG68K.C/TG68K_ALU.vhd:226:17  */
  assign n9629_o = n9553_o ? n9557_o : n9628_o;
  assign n9630_o = n9629_o[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:224:17  */
  assign n9631_o = n9549_o ? n9550_o : n9630_o;
  assign n9632_o = n9629_o[31:8];
  assign n9633_o = n9764_o[31:8];
  /* ../TG68K.C/TG68K_ALU.vhd:224:17  */
  assign n9634_o = n9549_o ? n9633_o : n9632_o;
  /* ../TG68K.C/TG68K_ALU.vhd:293:24  */
  assign n9639_o = exec[29];
  /* ../TG68K.C/TG68K_ALU.vhd:294:34  */
  assign n9640_o = sndopc[11];
  /* ../TG68K.C/TG68K_ALU.vhd:295:51  */
  assign n9641_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:295:62  */
  assign n9642_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:295:55  */
  assign n9643_o = {n9641_o, n9642_o};
  /* ../TG68K.C/TG68K_ALU.vhd:295:73  */
  assign n9644_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:295:66  */
  assign n9645_o = {n9643_o, n9644_o};
  /* ../TG68K.C/TG68K_ALU.vhd:295:84  */
  assign n9646_o = op1out[31:3];
  /* ../TG68K.C/TG68K_ALU.vhd:295:77  */
  assign n9647_o = {n9645_o, n9646_o};
  /* ../TG68K.C/TG68K_ALU.vhd:297:84  */
  assign n9648_o = sndopc[10:9];
  /* ../TG68K.C/TG68K_ALU.vhd:297:77  */
  assign n9650_o = {30'b000000000000000000000000000000, n9648_o};
  /* ../TG68K.C/TG68K_ALU.vhd:294:25  */
  assign n9651_o = n9640_o ? n9647_o : n9650_o;
  /* ../TG68K.C/TG68K_ALU.vhd:293:17  */
  assign n9652_o = n9639_o ? n9651_o : op1out;
  /* ../TG68K.C/TG68K_ALU.vhd:301:24  */
  assign n9653_o = exec[48];
  /* ../TG68K.C/TG68K_ALU.vhd:301:17  */
  assign n9656_o = n9653_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:309:24  */
  assign n9658_o = exec[78];
  /* ../TG68K.C/TG68K_ALU.vhd:310:65  */
  assign n9659_o = op2out[7:4];
  /* ../TG68K.C/TG68K_ALU.vhd:310:57  */
  assign n9661_o = {4'b0000, n9659_o};
  /* ../TG68K.C/TG68K_ALU.vhd:310:78  */
  assign n9663_o = {n9661_o, 4'b0000};
  /* ../TG68K.C/TG68K_ALU.vhd:310:95  */
  assign n9664_o = op2out[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:310:87  */
  assign n9665_o = {n9663_o, n9664_o};
  /* ../TG68K.C/TG68K_ALU.vhd:311:30  */
  assign n9666_o = ~execopc;
  /* ../TG68K.C/TG68K_ALU.vhd:311:43  */
  assign n9667_o = exec[53];
  /* ../TG68K.C/TG68K_ALU.vhd:311:55  */
  assign n9668_o = ~n9667_o;
  /* ../TG68K.C/TG68K_ALU.vhd:311:35  */
  assign n9669_o = n9666_o & n9668_o;
  /* ../TG68K.C/TG68K_ALU.vhd:311:68  */
  assign n9670_o = exec[29];
  /* ../TG68K.C/TG68K_ALU.vhd:311:82  */
  assign n9671_o = ~n9670_o;
  /* ../TG68K.C/TG68K_ALU.vhd:311:60  */
  assign n9672_o = n9669_o & n9671_o;
  /* ../TG68K.C/TG68K_ALU.vhd:312:38  */
  assign n9673_o = ~long_start;
  /* ../TG68K.C/TG68K_ALU.vhd:312:59  */
  assign n9675_o = exe_datatype == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:312:43  */
  assign n9676_o = n9673_o & n9675_o;
  /* ../TG68K.C/TG68K_ALU.vhd:312:73  */
  assign n9677_o = exec[50];
  /* ../TG68K.C/TG68K_ALU.vhd:312:81  */
  assign n9678_o = ~n9677_o;
  /* ../TG68K.C/TG68K_ALU.vhd:312:65  */
  assign n9679_o = n9676_o & n9678_o;
  /* ../TG68K.C/TG68K_ALU.vhd:314:41  */
  assign n9680_o = ~long_start;
  /* ../TG68K.C/TG68K_ALU.vhd:314:62  */
  assign n9682_o = exe_datatype == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:314:46  */
  assign n9683_o = n9680_o & n9682_o;
  /* ../TG68K.C/TG68K_ALU.vhd:314:77  */
  assign n9684_o = exec[47];
  /* ../TG68K.C/TG68K_ALU.vhd:314:93  */
  assign n9685_o = exec[46];
  /* ../TG68K.C/TG68K_ALU.vhd:314:86  */
  assign n9686_o = n9684_o | n9685_o;
  /* ../TG68K.C/TG68K_ALU.vhd:314:103  */
  assign n9687_o = n9686_o | movem_presub;
  /* ../TG68K.C/TG68K_ALU.vhd:314:68  */
  assign n9688_o = n9683_o & n9687_o;
  /* ../TG68K.C/TG68K_ALU.vhd:315:40  */
  assign n9689_o = exec[69];
  /* ../TG68K.C/TG68K_ALU.vhd:315:33  */
  assign n9692_o = n9689_o ? 32'b00000000000000000000000000000110 : 32'b00000000000000000000000000000100;
  /* ../TG68K.C/TG68K_ALU.vhd:314:25  */
  assign n9694_o = n9688_o ? n9692_o : 32'b00000000000000000000000000000010;
  /* ../TG68K.C/TG68K_ALU.vhd:312:25  */
  assign n9696_o = n9679_o ? 32'b00000000000000000000000000000001 : n9694_o;
  /* ../TG68K.C/TG68K_ALU.vhd:324:33  */
  assign n9697_o = exec[28];
  /* ../TG68K.C/TG68K_ALU.vhd:324:59  */
  assign n9698_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:324:50  */
  assign n9699_o = n9697_o & n9698_o;
  /* ../TG68K.C/TG68K_ALU.vhd:324:75  */
  assign n9700_o = exec[31];
  /* ../TG68K.C/TG68K_ALU.vhd:324:68  */
  assign n9701_o = n9699_o | n9700_o;
  /* ../TG68K.C/TG68K_ALU.vhd:324:25  */
  assign n9703_o = n9701_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:327:41  */
  assign n9704_o = exec[56];
  /* ../TG68K.C/TG68K_ALU.vhd:311:17  */
  assign n9705_o = n9672_o ? n9696_o : op2out;
  /* ../TG68K.C/TG68K_ALU.vhd:311:17  */
  assign n9706_o = n9672_o ? n9656_o : n9704_o;
  /* ../TG68K.C/TG68K_ALU.vhd:311:17  */
  assign n9707_o = n9672_o ? 1'b0 : n9703_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1316:25  */
  assign n9708_o = n9705_o[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:309:17  */
  assign n9709_o = n9658_o ? n9665_o : n9708_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1285:17  */
  assign n9710_o = n9705_o[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1283:1  */
  assign n9711_o = op2out[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:309:17  */
  assign n9712_o = n9658_o ? n9711_o : n9710_o;
  /* ../TG68K.C/TG68K_ALU.vhd:309:17  */
  assign n9714_o = n9658_o ? n9656_o : n9706_o;
  /* ../TG68K.C/TG68K_ALU.vhd:309:17  */
  assign n9715_o = n9658_o ? 1'b0 : n9707_o;
  /* ../TG68K.C/TG68K_ALU.vhd:331:24  */
  assign n9716_o = exec[69];
  /* ../TG68K.C/TG68K_ALU.vhd:331:43  */
  assign n9717_o = n9716_o | check_aligned;
  /* ../TG68K.C/TG68K_ALU.vhd:332:36  */
  assign n9718_o = ~movem_presub;
  /* ../TG68K.C/TG68K_ALU.vhd:333:64  */
  assign n9719_o = ~long_start;
  /* ../TG68K.C/TG68K_ALU.vhd:333:48  */
  assign n9720_o = non_aligned & n9719_o;
  assign n9722_o = {n9712_o, n9709_o};
  /* ../TG68K.C/TG68K_ALU.vhd:333:25  */
  assign n9723_o = n9720_o ? 32'b00000000000000000000000000000000 : n9722_o;
  /* ../TG68K.C/TG68K_ALU.vhd:337:64  */
  assign n9724_o = ~long_start;
  /* ../TG68K.C/TG68K_ALU.vhd:337:48  */
  assign n9725_o = non_aligned & n9724_o;
  /* ../TG68K.C/TG68K_ALU.vhd:338:44  */
  assign n9727_o = exe_datatype == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:338:27  */
  assign n9730_o = n9727_o ? 32'b00000000000000000000000000001000 : 32'b00000000000000000000000000000100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1010:17  */
  assign n9731_o = {n9712_o, n9709_o};
  /* ../TG68K.C/TG68K_ALU.vhd:337:25  */
  assign n9732_o = n9725_o ? n9730_o : n9731_o;
  /* ../TG68K.C/TG68K_ALU.vhd:332:19  */
  assign n9733_o = n9718_o ? n9723_o : n9732_o;
  assign n9734_o = {n9712_o, n9709_o};
  /* ../TG68K.C/TG68K_ALU.vhd:331:17  */
  assign n9735_o = n9717_o ? n9733_o : n9734_o;
  /* ../TG68K.C/TG68K_ALU.vhd:347:28  */
  assign n9736_o = ~opaddsub;
  /* ../TG68K.C/TG68K_ALU.vhd:347:33  */
  assign n9737_o = n9736_o | long_start;
  /* ../TG68K.C/TG68K_ALU.vhd:348:43  */
  assign n9739_o = {1'b0, addsub_b};
  /* ../TG68K.C/TG68K_ALU.vhd:348:57  */
  assign n9740_o = c_in[0];
  /* ../TG68K.C/TG68K_ALU.vhd:348:52  */
  assign n9741_o = {n9739_o, n9740_o};
  /* ../TG68K.C/TG68K_ALU.vhd:350:48  */
  assign n9743_o = {1'b0, addsub_b};
  /* ../TG68K.C/TG68K_ALU.vhd:350:62  */
  assign n9744_o = c_in[0];
  /* ../TG68K.C/TG68K_ALU.vhd:350:57  */
  assign n9745_o = {n9743_o, n9744_o};
  /* ../TG68K.C/TG68K_ALU.vhd:350:40  */
  assign n9746_o = ~n9745_o;
  /* ../TG68K.C/TG68K_ALU.vhd:347:17  */
  assign n9747_o = n9737_o ? n9741_o : n9746_o;
  /* ../TG68K.C/TG68K_ALU.vhd:352:36  */
  assign n9749_o = {1'b0, addsub_a};
  /* ../TG68K.C/TG68K_ALU.vhd:352:57  */
  assign n9750_o = notaddsub_b[0];
  /* ../TG68K.C/TG68K_ALU.vhd:352:45  */
  assign n9751_o = {n9749_o, n9750_o};
  /* ../TG68K.C/TG68K_ALU.vhd:352:61  */
  assign n9752_o = n9751_o + notaddsub_b;
  /* ../TG68K.C/TG68K_ALU.vhd:353:38  */
  assign n9753_o = add_result[9];
  /* ../TG68K.C/TG68K_ALU.vhd:353:54  */
  assign n9754_o = addsub_a[8];
  /* ../TG68K.C/TG68K_ALU.vhd:353:42  */
  assign n9755_o = n9753_o ^ n9754_o;
  /* ../TG68K.C/TG68K_ALU.vhd:353:70  */
  assign n9756_o = addsub_b[8];
  /* ../TG68K.C/TG68K_ALU.vhd:353:58  */
  assign n9757_o = n9755_o ^ n9756_o;
  /* ../TG68K.C/TG68K_ALU.vhd:354:38  */
  assign n9758_o = add_result[17];
  /* ../TG68K.C/TG68K_ALU.vhd:354:55  */
  assign n9759_o = addsub_a[16];
  /* ../TG68K.C/TG68K_ALU.vhd:354:43  */
  assign n9760_o = n9758_o ^ n9759_o;
  /* ../TG68K.C/TG68K_ALU.vhd:354:72  */
  assign n9761_o = addsub_b[16];
  /* ../TG68K.C/TG68K_ALU.vhd:354:60  */
  assign n9762_o = n9760_o ^ n9761_o;
  /* ../TG68K.C/TG68K_ALU.vhd:355:38  */
  assign n9763_o = add_result[33];
  /* ../TG68K.C/TG68K_ALU.vhd:356:39  */
  assign n9764_o = add_result[32:1];
  /* ../TG68K.C/TG68K_ALU.vhd:357:39  */
  assign n9765_o = c_in[1];
  /* ../TG68K.C/TG68K_ALU.vhd:357:57  */
  assign n9766_o = add_result[8];
  /* ../TG68K.C/TG68K_ALU.vhd:357:43  */
  assign n9767_o = n9765_o ^ n9766_o;
  /* ../TG68K.C/TG68K_ALU.vhd:357:73  */
  assign n9768_o = addsub_a[7];
  /* ../TG68K.C/TG68K_ALU.vhd:357:61  */
  assign n9769_o = n9767_o ^ n9768_o;
  /* ../TG68K.C/TG68K_ALU.vhd:357:89  */
  assign n9770_o = addsub_b[7];
  /* ../TG68K.C/TG68K_ALU.vhd:357:77  */
  assign n9771_o = n9769_o ^ n9770_o;
  /* ../TG68K.C/TG68K_ALU.vhd:358:39  */
  assign n9772_o = c_in[2];
  /* ../TG68K.C/TG68K_ALU.vhd:358:57  */
  assign n9773_o = add_result[16];
  /* ../TG68K.C/TG68K_ALU.vhd:358:43  */
  assign n9774_o = n9772_o ^ n9773_o;
  /* ../TG68K.C/TG68K_ALU.vhd:358:74  */
  assign n9775_o = addsub_a[15];
  /* ../TG68K.C/TG68K_ALU.vhd:358:62  */
  assign n9776_o = n9774_o ^ n9775_o;
  /* ../TG68K.C/TG68K_ALU.vhd:358:91  */
  assign n9777_o = addsub_b[15];
  /* ../TG68K.C/TG68K_ALU.vhd:358:79  */
  assign n9778_o = n9776_o ^ n9777_o;
  /* ../TG68K.C/TG68K_ALU.vhd:359:39  */
  assign n9779_o = c_in[3];
  /* ../TG68K.C/TG68K_ALU.vhd:359:57  */
  assign n9780_o = add_result[32];
  /* ../TG68K.C/TG68K_ALU.vhd:359:43  */
  assign n9781_o = n9779_o ^ n9780_o;
  /* ../TG68K.C/TG68K_ALU.vhd:359:74  */
  assign n9782_o = addsub_a[31];
  /* ../TG68K.C/TG68K_ALU.vhd:359:62  */
  assign n9783_o = n9781_o ^ n9782_o;
  /* ../TG68K.C/TG68K_ALU.vhd:359:91  */
  assign n9784_o = addsub_b[31];
  /* ../TG68K.C/TG68K_ALU.vhd:359:79  */
  assign n9785_o = n9783_o ^ n9784_o;
  /* ../TG68K.C/TG68K_ALU.vhd:360:30  */
  assign n9786_o = c_in[3:1];
  /* ../TG68K.C/TG68K_ALU.vhd:370:32  */
  assign n9790_o = c_in[1];
  /* ../TG68K.C/TG68K_ALU.vhd:370:46  */
  assign n9791_o = add_result[8:0];
  /* ../TG68K.C/TG68K_ALU.vhd:370:35  */
  assign n9792_o = {n9790_o, n9791_o};
  /* ../TG68K.C/TG68K_ALU.vhd:372:38  */
  assign n9793_o = op1out[4];
  /* ../TG68K.C/TG68K_ALU.vhd:372:52  */
  assign n9794_o = op2out[4];
  /* ../TG68K.C/TG68K_ALU.vhd:372:42  */
  assign n9795_o = n9793_o ^ n9794_o;
  /* ../TG68K.C/TG68K_ALU.vhd:372:67  */
  assign n9796_o = bcd_pur[5];
  /* ../TG68K.C/TG68K_ALU.vhd:372:56  */
  assign n9797_o = n9795_o ^ n9796_o;
  /* ../TG68K.C/TG68K_ALU.vhd:373:17  */
  assign n9800_o = halve_carry ? 4'b0110 : 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:376:27  */
  assign n9803_o = bcd_pur[9];
  assign n9805_o = n9801_o[7:4];
  /* ../TG68K.C/TG68K_ALU.vhd:376:17  */
  assign n9806_o = n9803_o ? 4'b0110 : n9805_o;
  assign n9807_o = n9801_o[8];
  /* ../TG68K.C/TG68K_ALU.vhd:379:24  */
  assign n9808_o = exec[12];
  /* ../TG68K.C/TG68K_ALU.vhd:380:47  */
  assign n9809_o = bcd_pur[8];
  /* ../TG68K.C/TG68K_ALU.vhd:380:36  */
  assign n9810_o = ~n9809_o;
  /* ../TG68K.C/TG68K_ALU.vhd:380:60  */
  assign n9811_o = bcd_a[7];
  /* ../TG68K.C/TG68K_ALU.vhd:380:51  */
  assign n9812_o = n9810_o & n9811_o;
  /* ../TG68K.C/TG68K_ALU.vhd:382:41  */
  assign n9813_o = bcd_pur[9:1];
  /* ../TG68K.C/TG68K_ALU.vhd:382:54  */
  assign n9814_o = n9813_o + bcd_kor;
  /* ../TG68K.C/TG68K_ALU.vhd:383:36  */
  assign n9815_o = bcd_pur[4];
  /* ../TG68K.C/TG68K_ALU.vhd:383:52  */
  assign n9816_o = bcd_pur[3];
  /* ../TG68K.C/TG68K_ALU.vhd:383:66  */
  assign n9817_o = bcd_pur[2];
  /* ../TG68K.C/TG68K_ALU.vhd:383:56  */
  assign n9818_o = n9816_o | n9817_o;
  /* ../TG68K.C/TG68K_ALU.vhd:383:40  */
  assign n9819_o = n9815_o & n9818_o;
  /* ../TG68K.C/TG68K_ALU.vhd:383:25  */
  assign n9821_o = n9819_o ? 4'b0110 : n9800_o;
  /* ../TG68K.C/TG68K_ALU.vhd:386:36  */
  assign n9822_o = bcd_pur[8];
  /* ../TG68K.C/TG68K_ALU.vhd:386:52  */
  assign n9823_o = bcd_pur[7];
  /* ../TG68K.C/TG68K_ALU.vhd:386:66  */
  assign n9824_o = bcd_pur[6];
  /* ../TG68K.C/TG68K_ALU.vhd:386:56  */
  assign n9825_o = n9823_o | n9824_o;
  /* ../TG68K.C/TG68K_ALU.vhd:386:81  */
  assign n9826_o = bcd_pur[5];
  /* ../TG68K.C/TG68K_ALU.vhd:386:96  */
  assign n9827_o = bcd_pur[4];
  /* ../TG68K.C/TG68K_ALU.vhd:386:85  */
  assign n9828_o = n9826_o & n9827_o;
  /* ../TG68K.C/TG68K_ALU.vhd:386:112  */
  assign n9829_o = bcd_pur[3];
  /* ../TG68K.C/TG68K_ALU.vhd:386:126  */
  assign n9830_o = bcd_pur[2];
  /* ../TG68K.C/TG68K_ALU.vhd:386:116  */
  assign n9831_o = n9829_o | n9830_o;
  /* ../TG68K.C/TG68K_ALU.vhd:386:100  */
  assign n9832_o = n9828_o & n9831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:386:70  */
  assign n9833_o = n9825_o | n9832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:386:40  */
  assign n9834_o = n9822_o & n9833_o;
  /* ../TG68K.C/TG68K_ALU.vhd:386:25  */
  assign n9836_o = n9834_o ? 4'b0110 : n9806_o;
  /* ../TG68K.C/TG68K_ALU.vhd:390:43  */
  assign n9837_o = bcd_pur[8];
  /* ../TG68K.C/TG68K_ALU.vhd:390:60  */
  assign n9838_o = bcd_a[7];
  /* ../TG68K.C/TG68K_ALU.vhd:390:51  */
  assign n9839_o = ~n9838_o;
  /* ../TG68K.C/TG68K_ALU.vhd:390:47  */
  assign n9840_o = n9837_o & n9839_o;
  /* ../TG68K.C/TG68K_ALU.vhd:392:41  */
  assign n9841_o = bcd_pur[9:1];
  /* ../TG68K.C/TG68K_ALU.vhd:392:54  */
  assign n9842_o = n9841_o - bcd_kor;
  assign n9843_o = {n9836_o, n9821_o};
  assign n9844_o = {n9806_o, n9800_o};
  /* ../TG68K.C/TG68K_ALU.vhd:379:17  */
  assign n9845_o = n9808_o ? n9843_o : n9844_o;
  /* ../TG68K.C/TG68K_ALU.vhd:379:17  */
  assign n9846_o = n9808_o ? n9812_o : n9840_o;
  /* ../TG68K.C/TG68K_ALU.vhd:379:17  */
  assign n9847_o = n9808_o ? n9814_o : n9842_o;
  /* ../TG68K.C/TG68K_ALU.vhd:394:23  */
  assign n9848_o = cpu[1];
  /* ../TG68K.C/TG68K_ALU.vhd:394:17  */
  assign n9850_o = n9848_o ? 1'b0 : n9846_o;
  /* ../TG68K.C/TG68K_ALU.vhd:397:39  */
  assign n9851_o = bcd_pur[9];
  /* ../TG68K.C/TG68K_ALU.vhd:397:51  */
  assign n9852_o = bcd_a[8];
  /* ../TG68K.C/TG68K_ALU.vhd:397:43  */
  assign n9853_o = n9851_o | n9852_o;
  /* ../TG68K.C/TG68K_ALU.vhd:409:44  */
  assign n9858_o = opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:410:41  */
  assign n9860_o = n9858_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:412:41  */
  assign n9862_o = n9858_o == 2'b11;
  assign n9863_o = {n9862_o, n9860_o};
  /* ../TG68K.C/TG68K_ALU.vhd:409:33  */
  always @*
    case (n9863_o)
      2'b10: n9866_o = 1'b0;
      2'b01: n9866_o = 1'b1;
      default: n9866_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:409:33  */
  always @*
    case (n9863_o)
      2'b10: n9870_o = 1'b1;
      2'b01: n9870_o = 1'b0;
      default: n9870_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:419:30  */
  assign n9876_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:419:33  */
  assign n9877_o = ~n9876_o;
  /* ../TG68K.C/TG68K_ALU.vhd:420:38  */
  assign n9878_o = exe_opcode[5:4];
  /* ../TG68K.C/TG68K_ALU.vhd:420:50  */
  assign n9880_o = n9878_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:421:53  */
  assign n9881_o = sndopc[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:423:58  */
  assign n9882_o = sndopc[2:0];
  /* ../TG68K.C/TG68K_ALU.vhd:423:51  */
  assign n9884_o = {2'b00, n9882_o};
  /* ../TG68K.C/TG68K_ALU.vhd:420:25  */
  assign n9885_o = n9880_o ? n9881_o : n9884_o;
  /* ../TG68K.C/TG68K_ALU.vhd:426:38  */
  assign n9886_o = exe_opcode[5:4];
  /* ../TG68K.C/TG68K_ALU.vhd:426:50  */
  assign n9888_o = n9886_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:427:53  */
  assign n9889_o = reg_qb[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:429:58  */
  assign n9890_o = reg_qb[2:0];
  /* ../TG68K.C/TG68K_ALU.vhd:429:51  */
  assign n9892_o = {2'b00, n9890_o};
  /* ../TG68K.C/TG68K_ALU.vhd:426:25  */
  assign n9893_o = n9888_o ? n9889_o : n9892_o;
  /* ../TG68K.C/TG68K_ALU.vhd:419:17  */
  assign n9894_o = n9877_o ? n9885_o : n9893_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:65  */
  assign n9900_o = ~one_bit_in;
  /* ../TG68K.C/TG68K_ALU.vhd:435:61  */
  assign n9901_o = bchg & n9900_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:81  */
  assign n9902_o = n9901_o | bset;
  /* ../TG68K.C/TG68K_ALU.vhd:456:42  */
  assign n9908_o = opcode[5:4];
  /* ../TG68K.C/TG68K_ALU.vhd:456:55  */
  assign n9910_o = n9908_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:456:33  */
  assign n9913_o = n9910_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:459:44  */
  assign n9915_o = opcode[10:8];
  /* ../TG68K.C/TG68K_ALU.vhd:460:41  */
  assign n9917_o = n9915_o == 3'b010;
  /* ../TG68K.C/TG68K_ALU.vhd:461:41  */
  assign n9919_o = n9915_o == 3'b011;
  /* ../TG68K.C/TG68K_ALU.vhd:463:41  */
  assign n9921_o = n9915_o == 3'b101;
  /* ../TG68K.C/TG68K_ALU.vhd:464:41  */
  assign n9923_o = n9915_o == 3'b110;
  /* ../TG68K.C/TG68K_ALU.vhd:465:41  */
  assign n9925_o = n9915_o == 3'b111;
  assign n9926_o = {n9925_o, n9923_o, n9921_o, n9919_o, n9917_o};
  /* ../TG68K.C/TG68K_ALU.vhd:459:33  */
  always @*
    case (n9926_o)
      5'b10000: n9929_o = 1'b0;
      5'b01000: n9929_o = 1'b1;
      5'b00100: n9929_o = 1'b0;
      5'b00010: n9929_o = 1'b0;
      5'b00001: n9929_o = 1'b0;
      default: n9929_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:459:33  */
  always @*
    case (n9926_o)
      5'b10000: n9933_o = 1'b0;
      5'b01000: n9933_o = 1'b0;
      5'b00100: n9933_o = 1'b0;
      5'b00010: n9933_o = 1'b0;
      5'b00001: n9933_o = 1'b1;
      default: n9933_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:459:33  */
  always @*
    case (n9926_o)
      5'b10000: n9937_o = 1'b1;
      5'b01000: n9937_o = 1'b0;
      5'b00100: n9937_o = 1'b0;
      5'b00010: n9937_o = 1'b0;
      5'b00001: n9937_o = 1'b0;
      default: n9937_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:459:33  */
  always @*
    case (n9926_o)
      5'b10000: n9941_o = 1'b0;
      5'b01000: n9941_o = 1'b0;
      5'b00100: n9941_o = 1'b0;
      5'b00010: n9941_o = 1'b1;
      5'b00001: n9941_o = 1'b0;
      default: n9941_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:459:33  */
  always @*
    case (n9926_o)
      5'b10000: n9945_o = 1'b0;
      5'b01000: n9945_o = 1'b0;
      5'b00100: n9945_o = 1'b1;
      5'b00010: n9945_o = 1'b0;
      5'b00001: n9945_o = 1'b0;
      default: n9945_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:459:33  */
  always @*
    case (n9926_o)
      5'b10000: n9948_o = 1'b1;
      5'b01000: n9948_o = n9913_o;
      5'b00100: n9948_o = n9913_o;
      5'b00010: n9948_o = n9913_o;
      5'b00001: n9948_o = n9913_o;
      default: n9948_o = n9913_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:469:42  */
  assign n9949_o = opcode[4:3];
  /* ../TG68K.C/TG68K_ALU.vhd:469:54  */
  assign n9951_o = n9949_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:469:33  */
  assign n9954_o = n9951_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:472:53  */
  assign n9956_o = result[39:32];
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n9974_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n9976_o = $unsigned(5'b00000) > $unsigned(n9974_o);
  assign n9979_o = reg_qb[0];
  assign n9980_o = bf_set2[0];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n9981_o = bf_ins ? n9979_o : n9980_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n9982_o = n9976_o ? 1'b0 : n9981_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n9987_o = n9976_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n9990_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n9992_o = $unsigned(5'b00001) > $unsigned(n9990_o);
  assign n9995_o = reg_qb[1];
  assign n9996_o = bf_set2[1];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n9997_o = bf_ins ? n9995_o : n9996_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n9998_o = n9992_o ? 1'b0 : n9997_o;
  assign n10002_o = n9988_o[1];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10003_o = n9992_o ? 1'b1 : n10002_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10005_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10007_o = $unsigned(5'b00010) > $unsigned(n10005_o);
  assign n10010_o = reg_qb[2];
  assign n10011_o = bf_set2[2];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10012_o = bf_ins ? n10010_o : n10011_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10013_o = n10007_o ? 1'b0 : n10012_o;
  assign n10017_o = n9988_o[2];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10018_o = n10007_o ? 1'b1 : n10017_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10020_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10022_o = $unsigned(5'b00011) > $unsigned(n10020_o);
  assign n10025_o = reg_qb[3];
  assign n10026_o = bf_set2[3];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10027_o = bf_ins ? n10025_o : n10026_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10028_o = n10022_o ? 1'b0 : n10027_o;
  assign n10032_o = n9988_o[3];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10033_o = n10022_o ? 1'b1 : n10032_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10035_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10037_o = $unsigned(5'b00100) > $unsigned(n10035_o);
  assign n10040_o = reg_qb[4];
  assign n10041_o = bf_set2[4];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10042_o = bf_ins ? n10040_o : n10041_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10043_o = n10037_o ? 1'b0 : n10042_o;
  assign n10047_o = n9988_o[4];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10048_o = n10037_o ? 1'b1 : n10047_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10050_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10052_o = $unsigned(5'b00101) > $unsigned(n10050_o);
  assign n10055_o = reg_qb[5];
  assign n10056_o = bf_set2[5];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10057_o = bf_ins ? n10055_o : n10056_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10058_o = n10052_o ? 1'b0 : n10057_o;
  assign n10062_o = n9988_o[5];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10063_o = n10052_o ? 1'b1 : n10062_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10065_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10067_o = $unsigned(5'b00110) > $unsigned(n10065_o);
  assign n10070_o = reg_qb[6];
  assign n10071_o = bf_set2[6];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10072_o = bf_ins ? n10070_o : n10071_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10073_o = n10067_o ? 1'b0 : n10072_o;
  assign n10077_o = n9988_o[6];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10078_o = n10067_o ? 1'b1 : n10077_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10080_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10082_o = $unsigned(5'b00111) > $unsigned(n10080_o);
  assign n10085_o = reg_qb[7];
  assign n10086_o = bf_set2[7];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10087_o = bf_ins ? n10085_o : n10086_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10088_o = n10082_o ? 1'b0 : n10087_o;
  assign n10092_o = n9988_o[7];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10093_o = n10082_o ? 1'b1 : n10092_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10095_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10097_o = $unsigned(5'b01000) > $unsigned(n10095_o);
  assign n10100_o = reg_qb[8];
  assign n10101_o = bf_set2[8];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10102_o = bf_ins ? n10100_o : n10101_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10103_o = n10097_o ? 1'b0 : n10102_o;
  assign n10107_o = n9988_o[8];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10108_o = n10097_o ? 1'b1 : n10107_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10110_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10112_o = $unsigned(5'b01001) > $unsigned(n10110_o);
  assign n10115_o = reg_qb[9];
  assign n10116_o = bf_set2[9];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10117_o = bf_ins ? n10115_o : n10116_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10118_o = n10112_o ? 1'b0 : n10117_o;
  assign n10122_o = n9988_o[9];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10123_o = n10112_o ? 1'b1 : n10122_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10125_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10127_o = $unsigned(5'b01010) > $unsigned(n10125_o);
  assign n10130_o = reg_qb[10];
  assign n10131_o = bf_set2[10];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10132_o = bf_ins ? n10130_o : n10131_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10133_o = n10127_o ? 1'b0 : n10132_o;
  assign n10137_o = n9988_o[10];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10138_o = n10127_o ? 1'b1 : n10137_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10140_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10142_o = $unsigned(5'b01011) > $unsigned(n10140_o);
  assign n10145_o = reg_qb[11];
  assign n10146_o = bf_set2[11];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10147_o = bf_ins ? n10145_o : n10146_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10148_o = n10142_o ? 1'b0 : n10147_o;
  assign n10152_o = n9988_o[11];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10153_o = n10142_o ? 1'b1 : n10152_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10155_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10157_o = $unsigned(5'b01100) > $unsigned(n10155_o);
  assign n10160_o = reg_qb[12];
  assign n10161_o = bf_set2[12];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10162_o = bf_ins ? n10160_o : n10161_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10163_o = n10157_o ? 1'b0 : n10162_o;
  assign n10167_o = n9988_o[12];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10168_o = n10157_o ? 1'b1 : n10167_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10170_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10172_o = $unsigned(5'b01101) > $unsigned(n10170_o);
  assign n10175_o = reg_qb[13];
  assign n10176_o = bf_set2[13];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10177_o = bf_ins ? n10175_o : n10176_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10178_o = n10172_o ? 1'b0 : n10177_o;
  assign n10182_o = n9988_o[13];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10183_o = n10172_o ? 1'b1 : n10182_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10185_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10187_o = $unsigned(5'b01110) > $unsigned(n10185_o);
  assign n10190_o = reg_qb[14];
  assign n10191_o = bf_set2[14];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10192_o = bf_ins ? n10190_o : n10191_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10193_o = n10187_o ? 1'b0 : n10192_o;
  assign n10197_o = n9988_o[14];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10198_o = n10187_o ? 1'b1 : n10197_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10200_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10202_o = $unsigned(5'b01111) > $unsigned(n10200_o);
  assign n10205_o = reg_qb[15];
  assign n10206_o = bf_set2[15];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10207_o = bf_ins ? n10205_o : n10206_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10208_o = n10202_o ? 1'b0 : n10207_o;
  assign n10212_o = n9988_o[15];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10213_o = n10202_o ? 1'b1 : n10212_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10215_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10217_o = $unsigned(5'b10000) > $unsigned(n10215_o);
  assign n10220_o = reg_qb[16];
  assign n10221_o = bf_set2[16];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10222_o = bf_ins ? n10220_o : n10221_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10223_o = n10217_o ? 1'b0 : n10222_o;
  assign n10227_o = n9988_o[16];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10228_o = n10217_o ? 1'b1 : n10227_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10230_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10232_o = $unsigned(5'b10001) > $unsigned(n10230_o);
  assign n10235_o = reg_qb[17];
  assign n10236_o = bf_set2[17];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10237_o = bf_ins ? n10235_o : n10236_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10238_o = n10232_o ? 1'b0 : n10237_o;
  assign n10242_o = n9988_o[17];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10243_o = n10232_o ? 1'b1 : n10242_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10245_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10247_o = $unsigned(5'b10010) > $unsigned(n10245_o);
  assign n10250_o = reg_qb[18];
  assign n10251_o = bf_set2[18];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10252_o = bf_ins ? n10250_o : n10251_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10253_o = n10247_o ? 1'b0 : n10252_o;
  assign n10257_o = n9988_o[18];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10258_o = n10247_o ? 1'b1 : n10257_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10260_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10262_o = $unsigned(5'b10011) > $unsigned(n10260_o);
  assign n10265_o = reg_qb[19];
  assign n10266_o = bf_set2[19];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10267_o = bf_ins ? n10265_o : n10266_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10268_o = n10262_o ? 1'b0 : n10267_o;
  assign n10272_o = n9988_o[19];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10273_o = n10262_o ? 1'b1 : n10272_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10275_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10277_o = $unsigned(5'b10100) > $unsigned(n10275_o);
  assign n10280_o = reg_qb[20];
  assign n10281_o = bf_set2[20];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10282_o = bf_ins ? n10280_o : n10281_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10283_o = n10277_o ? 1'b0 : n10282_o;
  assign n10287_o = n9988_o[20];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10288_o = n10277_o ? 1'b1 : n10287_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10290_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10292_o = $unsigned(5'b10101) > $unsigned(n10290_o);
  assign n10295_o = reg_qb[21];
  assign n10296_o = bf_set2[21];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10297_o = bf_ins ? n10295_o : n10296_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10298_o = n10292_o ? 1'b0 : n10297_o;
  assign n10302_o = n9988_o[21];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10303_o = n10292_o ? 1'b1 : n10302_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10305_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10307_o = $unsigned(5'b10110) > $unsigned(n10305_o);
  assign n10310_o = reg_qb[22];
  assign n10311_o = bf_set2[22];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10312_o = bf_ins ? n10310_o : n10311_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10313_o = n10307_o ? 1'b0 : n10312_o;
  assign n10317_o = n9988_o[22];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10318_o = n10307_o ? 1'b1 : n10317_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10320_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10322_o = $unsigned(5'b10111) > $unsigned(n10320_o);
  assign n10325_o = reg_qb[23];
  assign n10326_o = bf_set2[23];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10327_o = bf_ins ? n10325_o : n10326_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10328_o = n10322_o ? 1'b0 : n10327_o;
  assign n10332_o = n9988_o[23];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10333_o = n10322_o ? 1'b1 : n10332_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10335_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10337_o = $unsigned(5'b11000) > $unsigned(n10335_o);
  assign n10340_o = reg_qb[24];
  assign n10341_o = bf_set2[24];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10342_o = bf_ins ? n10340_o : n10341_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10343_o = n10337_o ? 1'b0 : n10342_o;
  assign n10347_o = n9988_o[24];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10348_o = n10337_o ? 1'b1 : n10347_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10350_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10352_o = $unsigned(5'b11001) > $unsigned(n10350_o);
  assign n10355_o = reg_qb[25];
  assign n10356_o = bf_set2[25];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10357_o = bf_ins ? n10355_o : n10356_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10358_o = n10352_o ? 1'b0 : n10357_o;
  assign n10362_o = n9988_o[25];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10363_o = n10352_o ? 1'b1 : n10362_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10365_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10367_o = $unsigned(5'b11010) > $unsigned(n10365_o);
  assign n10370_o = reg_qb[26];
  assign n10371_o = bf_set2[26];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10372_o = bf_ins ? n10370_o : n10371_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10373_o = n10367_o ? 1'b0 : n10372_o;
  assign n10377_o = n9988_o[26];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10378_o = n10367_o ? 1'b1 : n10377_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10380_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10382_o = $unsigned(5'b11011) > $unsigned(n10380_o);
  assign n10385_o = reg_qb[27];
  assign n10386_o = bf_set2[27];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10387_o = bf_ins ? n10385_o : n10386_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10388_o = n10382_o ? 1'b0 : n10387_o;
  assign n10392_o = n9988_o[27];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10393_o = n10382_o ? 1'b1 : n10392_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10395_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10397_o = $unsigned(5'b11100) > $unsigned(n10395_o);
  assign n10400_o = reg_qb[28];
  assign n10401_o = bf_set2[28];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10402_o = bf_ins ? n10400_o : n10401_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10403_o = n10397_o ? 1'b0 : n10402_o;
  assign n10407_o = n9988_o[28];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10408_o = n10397_o ? 1'b1 : n10407_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10410_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10412_o = $unsigned(5'b11101) > $unsigned(n10410_o);
  assign n10415_o = reg_qb[29];
  assign n10416_o = bf_set2[29];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10417_o = bf_ins ? n10415_o : n10416_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10418_o = n10412_o ? 1'b0 : n10417_o;
  assign n10422_o = n9988_o[29];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10423_o = n10412_o ? 1'b1 : n10422_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10425_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10427_o = $unsigned(5'b11110) > $unsigned(n10425_o);
  assign n10430_o = reg_qb[30];
  assign n10431_o = bf_set2[30];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10432_o = bf_ins ? n10430_o : n10431_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10433_o = n10427_o ? 1'b0 : n10432_o;
  assign n10434_o = reg_qb[31];
  assign n10435_o = bf_set2[31];
  /* ../TG68K.C/TG68K_ALU.vhd:476:17  */
  assign n10436_o = bf_ins ? n10434_o : n10435_o;
  assign n10437_o = n9988_o[30];
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10438_o = n10427_o ? 1'b1 : n10437_o;
  assign n10439_o = n9988_o[31];
  /* ../TG68K.C/TG68K_ALU.vhd:490:38  */
  assign n10440_o = bf_width[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:490:29  */
  assign n10442_o = $unsigned(5'b11111) > $unsigned(n10440_o);
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10445_o = n10442_o ? 1'b0 : n10436_o;
  /* ../TG68K.C/TG68K_ALU.vhd:490:25  */
  assign n10446_o = n10442_o ? 1'b1 : n10439_o;
  /* ../TG68K.C/TG68K_ALU.vhd:496:37  */
  assign n10448_o = bf_width[4:0];  // trunc
  /* ../TG68K.C/TG68K_ALU.vhd:497:32  */
  assign n10451_o = bf_exts & bf_nflag;
  /* ../TG68K.C/TG68K_ALU.vhd:498:47  */
  assign n10452_o = datareg | unshifted_bitmask;
  /* ../TG68K.C/TG68K_ALU.vhd:497:17  */
  assign n10453_o = n10451_o ? n10452_o : datareg;
  /* ../TG68K.C/TG68K_ALU.vhd:504:30  */
  assign n10454_o = bf_loffset[4];
  /* ../TG68K.C/TG68K_ALU.vhd:505:57  */
  assign n10455_o = unshifted_bitmask[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:505:88  */
  assign n10456_o = unshifted_bitmask[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:505:70  */
  assign n10457_o = {n10455_o, n10456_o};
  /* ../TG68K.C/TG68K_ALU.vhd:504:17  */
  assign n10458_o = n10454_o ? n10457_o : unshifted_bitmask;
  /* ../TG68K.C/TG68K_ALU.vhd:509:30  */
  assign n10459_o = bf_loffset[3];
  /* ../TG68K.C/TG68K_ALU.vhd:510:64  */
  assign n10460_o = bitmaskmux3[23:0];
  /* ../TG68K.C/TG68K_ALU.vhd:510:89  */
  assign n10461_o = bitmaskmux3[31:24];
  /* ../TG68K.C/TG68K_ALU.vhd:510:77  */
  assign n10462_o = {n10460_o, n10461_o};
  /* ../TG68K.C/TG68K_ALU.vhd:509:17  */
  assign n10463_o = n10459_o ? n10462_o : bitmaskmux3;
  /* ../TG68K.C/TG68K_ALU.vhd:514:30  */
  assign n10464_o = bf_loffset[2];
  /* ../TG68K.C/TG68K_ALU.vhd:515:51  */
  assign n10466_o = {bitmaskmux2, 4'b1111};
  /* ../TG68K.C/TG68K_ALU.vhd:517:71  */
  assign n10467_o = bitmaskmux2[31:28];
  assign n10468_o = n10466_o[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:516:25  */
  assign n10469_o = bf_d32 ? n10467_o : n10468_o;
  assign n10470_o = n10466_o[35:4];
  /* ../TG68K.C/TG68K_ALU.vhd:520:46  */
  assign n10472_o = {4'b1111, bitmaskmux2};
  assign n10473_o = {n10470_o, n10469_o};
  /* ../TG68K.C/TG68K_ALU.vhd:514:17  */
  assign n10474_o = n10464_o ? n10473_o : n10472_o;
  /* ../TG68K.C/TG68K_ALU.vhd:522:30  */
  assign n10475_o = bf_loffset[1];
  /* ../TG68K.C/TG68K_ALU.vhd:523:51  */
  assign n10477_o = {bitmaskmux1, 2'b11};
  /* ../TG68K.C/TG68K_ALU.vhd:525:71  */
  assign n10478_o = bitmaskmux1[31:30];
  assign n10479_o = n10477_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:524:25  */
  assign n10480_o = bf_d32 ? n10478_o : n10479_o;
  assign n10481_o = n10477_o[37:2];
  /* ../TG68K.C/TG68K_ALU.vhd:528:44  */
  assign n10483_o = {2'b11, bitmaskmux1};
  assign n10484_o = {n10481_o, n10480_o};
  /* ../TG68K.C/TG68K_ALU.vhd:522:17  */
  assign n10485_o = n10475_o ? n10484_o : n10483_o;
  /* ../TG68K.C/TG68K_ALU.vhd:530:30  */
  assign n10486_o = bf_loffset[0];
  /* ../TG68K.C/TG68K_ALU.vhd:531:47  */
  assign n10488_o = {1'b1, bitmaskmux0};
  /* ../TG68K.C/TG68K_ALU.vhd:531:59  */
  assign n10490_o = {n10488_o, 1'b1};
  /* ../TG68K.C/TG68K_ALU.vhd:533:66  */
  assign n10491_o = bitmaskmux0[31];
  assign n10492_o = n10490_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:532:25  */
  assign n10493_o = bf_d32 ? n10491_o : n10492_o;
  assign n10494_o = n10490_o[39:1];
  /* ../TG68K.C/TG68K_ALU.vhd:536:48  */
  assign n10496_o = {2'b11, bitmaskmux0};
  assign n10497_o = {n10494_o, n10493_o};
  /* ../TG68K.C/TG68K_ALU.vhd:530:17  */
  assign n10498_o = n10486_o ? n10497_o : n10496_o;
  /* ../TG68K.C/TG68K_ALU.vhd:541:35  */
  assign n10499_o = {bf_ext_in, op2out};
  /* ../TG68K.C/TG68K_ALU.vhd:543:54  */
  assign n10500_o = op2out[7:0];
  assign n10501_o = n10499_o[39:32];
  /* ../TG68K.C/TG68K_ALU.vhd:542:17  */
  assign n10502_o = bf_s32 ? n10500_o : n10501_o;
  assign n10503_o = n10499_o[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:546:28  */
  assign n10504_o = bf_shift[0];
  /* ../TG68K.C/TG68K_ALU.vhd:547:40  */
  assign n10505_o = shift[0];
  /* ../TG68K.C/TG68K_ALU.vhd:547:49  */
  assign n10506_o = shift[39:1];
  /* ../TG68K.C/TG68K_ALU.vhd:547:43  */
  assign n10507_o = {n10505_o, n10506_o};
  /* ../TG68K.C/TG68K_ALU.vhd:546:17  */
  assign n10508_o = n10504_o ? n10507_o : shift;
  /* ../TG68K.C/TG68K_ALU.vhd:551:28  */
  assign n10509_o = bf_shift[1];
  /* ../TG68K.C/TG68K_ALU.vhd:552:41  */
  assign n10510_o = inmux0[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:552:60  */
  assign n10511_o = inmux0[39:2];
  /* ../TG68K.C/TG68K_ALU.vhd:552:53  */
  assign n10512_o = {n10510_o, n10511_o};
  /* ../TG68K.C/TG68K_ALU.vhd:551:17  */
  assign n10513_o = n10509_o ? n10512_o : inmux0;
  /* ../TG68K.C/TG68K_ALU.vhd:556:28  */
  assign n10514_o = bf_shift[2];
  /* ../TG68K.C/TG68K_ALU.vhd:557:41  */
  assign n10515_o = inmux1[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:557:60  */
  assign n10516_o = inmux1[39:4];
  /* ../TG68K.C/TG68K_ALU.vhd:557:53  */
  assign n10517_o = {n10515_o, n10516_o};
  /* ../TG68K.C/TG68K_ALU.vhd:556:17  */
  assign n10518_o = n10514_o ? n10517_o : inmux1;
  /* ../TG68K.C/TG68K_ALU.vhd:561:28  */
  assign n10519_o = bf_shift[3];
  /* ../TG68K.C/TG68K_ALU.vhd:562:41  */
  assign n10520_o = inmux2[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:562:60  */
  assign n10521_o = inmux2[31:8];
  /* ../TG68K.C/TG68K_ALU.vhd:562:53  */
  assign n10522_o = {n10520_o, n10521_o};
  /* ../TG68K.C/TG68K_ALU.vhd:564:41  */
  assign n10523_o = inmux2[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:561:17  */
  assign n10524_o = n10519_o ? n10522_o : n10523_o;
  /* ../TG68K.C/TG68K_ALU.vhd:566:28  */
  assign n10525_o = bf_shift[4];
  /* ../TG68K.C/TG68K_ALU.vhd:567:55  */
  assign n10526_o = inmux3[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:567:75  */
  assign n10527_o = inmux3[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:567:68  */
  assign n10528_o = {n10526_o, n10527_o};
  /* ../TG68K.C/TG68K_ALU.vhd:566:17  */
  assign n10529_o = n10525_o ? n10528_o : inmux3;
  /* ../TG68K.C/TG68K_ALU.vhd:574:56  */
  assign n10530_o = bf_set2[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:576:48  */
  assign n10531_o = ~op2out;
  /* ../TG68K.C/TG68K_ALU.vhd:577:49  */
  assign n10532_o = ~bf_ext_in;
  assign n10533_o = {n10532_o, n10531_o};
  assign n10536_o = {n10530_o, bf_set2};
  /* ../TG68K.C/TG68K_ALU.vhd:586:48  */
  assign n10540_o = {bf_ext_in, op1out};
  /* ../TG68K.C/TG68K_ALU.vhd:588:48  */
  assign n10541_o = {bf_ext_in, op2out};
  /* ../TG68K.C/TG68K_ALU.vhd:585:17  */
  assign n10542_o = bf_ins ? n10540_o : n10541_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10543_o = shifted_bitmask[0];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10544_o = result_tmp[0];
  assign n10545_o = n10538_o[0];
  assign n10546_o = n10536_o[0];
  assign n10547_o = n10533_o[0];
  assign n10548_o = n10534_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10549_o = bf_bchg ? n10547_o : n10548_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10550_o = bf_ins ? n10546_o : n10549_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10551_o = bf_bset ? n10545_o : n10550_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10552_o = n10543_o ? n10544_o : n10551_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10560_o = shifted_bitmask[1];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10561_o = result_tmp[1];
  assign n10562_o = n10538_o[1];
  assign n10563_o = n10536_o[1];
  assign n10564_o = n10533_o[1];
  assign n10565_o = n10534_o[1];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10566_o = bf_bchg ? n10564_o : n10565_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10567_o = bf_ins ? n10563_o : n10566_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10568_o = bf_bset ? n10562_o : n10567_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10569_o = n10560_o ? n10561_o : n10568_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10577_o = shifted_bitmask[2];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10578_o = result_tmp[2];
  assign n10579_o = n10538_o[2];
  assign n10580_o = n10536_o[2];
  assign n10581_o = n10533_o[2];
  assign n10582_o = n10534_o[2];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10583_o = bf_bchg ? n10581_o : n10582_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10584_o = bf_ins ? n10580_o : n10583_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10585_o = bf_bset ? n10579_o : n10584_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10586_o = n10577_o ? n10578_o : n10585_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10594_o = shifted_bitmask[3];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10595_o = result_tmp[3];
  assign n10596_o = n10538_o[3];
  assign n10597_o = n10536_o[3];
  assign n10598_o = n10533_o[3];
  assign n10599_o = n10534_o[3];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10600_o = bf_bchg ? n10598_o : n10599_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10601_o = bf_ins ? n10597_o : n10600_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10602_o = bf_bset ? n10596_o : n10601_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10603_o = n10594_o ? n10595_o : n10602_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10611_o = shifted_bitmask[4];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10612_o = result_tmp[4];
  assign n10613_o = n10538_o[4];
  assign n10614_o = n10536_o[4];
  assign n10615_o = n10533_o[4];
  assign n10616_o = n10534_o[4];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10617_o = bf_bchg ? n10615_o : n10616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10618_o = bf_ins ? n10614_o : n10617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10619_o = bf_bset ? n10613_o : n10618_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10620_o = n10611_o ? n10612_o : n10619_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10628_o = shifted_bitmask[5];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10629_o = result_tmp[5];
  assign n10630_o = n10538_o[5];
  assign n10631_o = n10536_o[5];
  assign n10632_o = n10533_o[5];
  assign n10633_o = n10534_o[5];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10634_o = bf_bchg ? n10632_o : n10633_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10635_o = bf_ins ? n10631_o : n10634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10636_o = bf_bset ? n10630_o : n10635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10637_o = n10628_o ? n10629_o : n10636_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10645_o = shifted_bitmask[6];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10646_o = result_tmp[6];
  assign n10647_o = n10538_o[6];
  assign n10648_o = n10536_o[6];
  assign n10649_o = n10533_o[6];
  assign n10650_o = n10534_o[6];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10651_o = bf_bchg ? n10649_o : n10650_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10652_o = bf_ins ? n10648_o : n10651_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10653_o = bf_bset ? n10647_o : n10652_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10654_o = n10645_o ? n10646_o : n10653_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10662_o = shifted_bitmask[7];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10663_o = result_tmp[7];
  assign n10664_o = n10538_o[7];
  assign n10665_o = n10536_o[7];
  assign n10666_o = n10533_o[7];
  assign n10667_o = n10534_o[7];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10668_o = bf_bchg ? n10666_o : n10667_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10669_o = bf_ins ? n10665_o : n10668_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10670_o = bf_bset ? n10664_o : n10669_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10671_o = n10662_o ? n10663_o : n10670_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10679_o = shifted_bitmask[8];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10680_o = result_tmp[8];
  assign n10681_o = n10538_o[8];
  assign n10682_o = n10536_o[8];
  assign n10683_o = n10533_o[8];
  assign n10684_o = n10534_o[8];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10685_o = bf_bchg ? n10683_o : n10684_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10686_o = bf_ins ? n10682_o : n10685_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10687_o = bf_bset ? n10681_o : n10686_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10688_o = n10679_o ? n10680_o : n10687_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10696_o = shifted_bitmask[9];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10697_o = result_tmp[9];
  assign n10698_o = n10538_o[9];
  assign n10699_o = n10536_o[9];
  assign n10700_o = n10533_o[9];
  assign n10701_o = n10534_o[9];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10702_o = bf_bchg ? n10700_o : n10701_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10703_o = bf_ins ? n10699_o : n10702_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10704_o = bf_bset ? n10698_o : n10703_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10705_o = n10696_o ? n10697_o : n10704_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10713_o = shifted_bitmask[10];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10714_o = result_tmp[10];
  assign n10715_o = n10538_o[10];
  assign n10716_o = n10536_o[10];
  assign n10717_o = n10533_o[10];
  assign n10718_o = n10534_o[10];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10719_o = bf_bchg ? n10717_o : n10718_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10720_o = bf_ins ? n10716_o : n10719_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10721_o = bf_bset ? n10715_o : n10720_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10722_o = n10713_o ? n10714_o : n10721_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10730_o = shifted_bitmask[11];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10731_o = result_tmp[11];
  assign n10732_o = n10538_o[11];
  assign n10733_o = n10536_o[11];
  assign n10734_o = n10533_o[11];
  assign n10735_o = n10534_o[11];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10736_o = bf_bchg ? n10734_o : n10735_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10737_o = bf_ins ? n10733_o : n10736_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10738_o = bf_bset ? n10732_o : n10737_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10739_o = n10730_o ? n10731_o : n10738_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10747_o = shifted_bitmask[12];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10748_o = result_tmp[12];
  assign n10749_o = n10538_o[12];
  assign n10750_o = n10536_o[12];
  assign n10751_o = n10533_o[12];
  assign n10752_o = n10534_o[12];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10753_o = bf_bchg ? n10751_o : n10752_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10754_o = bf_ins ? n10750_o : n10753_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10755_o = bf_bset ? n10749_o : n10754_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10756_o = n10747_o ? n10748_o : n10755_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10764_o = shifted_bitmask[13];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10765_o = result_tmp[13];
  assign n10766_o = n10538_o[13];
  assign n10767_o = n10536_o[13];
  assign n10768_o = n10533_o[13];
  assign n10769_o = n10534_o[13];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10770_o = bf_bchg ? n10768_o : n10769_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10771_o = bf_ins ? n10767_o : n10770_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10772_o = bf_bset ? n10766_o : n10771_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10773_o = n10764_o ? n10765_o : n10772_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10781_o = shifted_bitmask[14];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10782_o = result_tmp[14];
  assign n10783_o = n10538_o[14];
  assign n10784_o = n10536_o[14];
  assign n10785_o = n10533_o[14];
  assign n10786_o = n10534_o[14];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10787_o = bf_bchg ? n10785_o : n10786_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10788_o = bf_ins ? n10784_o : n10787_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10789_o = bf_bset ? n10783_o : n10788_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10790_o = n10781_o ? n10782_o : n10789_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10798_o = shifted_bitmask[15];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10799_o = result_tmp[15];
  assign n10800_o = n10538_o[15];
  assign n10801_o = n10536_o[15];
  assign n10802_o = n10533_o[15];
  assign n10803_o = n10534_o[15];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10804_o = bf_bchg ? n10802_o : n10803_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10805_o = bf_ins ? n10801_o : n10804_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10806_o = bf_bset ? n10800_o : n10805_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10807_o = n10798_o ? n10799_o : n10806_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10815_o = shifted_bitmask[16];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10816_o = result_tmp[16];
  assign n10817_o = n10538_o[16];
  assign n10818_o = n10536_o[16];
  assign n10819_o = n10533_o[16];
  assign n10820_o = n10534_o[16];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10821_o = bf_bchg ? n10819_o : n10820_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10822_o = bf_ins ? n10818_o : n10821_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10823_o = bf_bset ? n10817_o : n10822_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10824_o = n10815_o ? n10816_o : n10823_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10832_o = shifted_bitmask[17];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10833_o = result_tmp[17];
  assign n10834_o = n10538_o[17];
  assign n10835_o = n10536_o[17];
  assign n10836_o = n10533_o[17];
  assign n10837_o = n10534_o[17];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10838_o = bf_bchg ? n10836_o : n10837_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10839_o = bf_ins ? n10835_o : n10838_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10840_o = bf_bset ? n10834_o : n10839_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10841_o = n10832_o ? n10833_o : n10840_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10849_o = shifted_bitmask[18];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10850_o = result_tmp[18];
  assign n10851_o = n10538_o[18];
  assign n10852_o = n10536_o[18];
  assign n10853_o = n10533_o[18];
  assign n10854_o = n10534_o[18];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10855_o = bf_bchg ? n10853_o : n10854_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10856_o = bf_ins ? n10852_o : n10855_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10857_o = bf_bset ? n10851_o : n10856_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10858_o = n10849_o ? n10850_o : n10857_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10866_o = shifted_bitmask[19];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10867_o = result_tmp[19];
  assign n10868_o = n10538_o[19];
  assign n10869_o = n10536_o[19];
  assign n10870_o = n10533_o[19];
  assign n10871_o = n10534_o[19];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10872_o = bf_bchg ? n10870_o : n10871_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10873_o = bf_ins ? n10869_o : n10872_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10874_o = bf_bset ? n10868_o : n10873_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10875_o = n10866_o ? n10867_o : n10874_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10883_o = shifted_bitmask[20];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10884_o = result_tmp[20];
  assign n10885_o = n10538_o[20];
  assign n10886_o = n10536_o[20];
  assign n10887_o = n10533_o[20];
  assign n10888_o = n10534_o[20];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10889_o = bf_bchg ? n10887_o : n10888_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10890_o = bf_ins ? n10886_o : n10889_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10891_o = bf_bset ? n10885_o : n10890_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10892_o = n10883_o ? n10884_o : n10891_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10900_o = shifted_bitmask[21];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10901_o = result_tmp[21];
  assign n10902_o = n10538_o[21];
  assign n10903_o = n10536_o[21];
  assign n10904_o = n10533_o[21];
  assign n10905_o = n10534_o[21];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10906_o = bf_bchg ? n10904_o : n10905_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10907_o = bf_ins ? n10903_o : n10906_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10908_o = bf_bset ? n10902_o : n10907_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10909_o = n10900_o ? n10901_o : n10908_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10917_o = shifted_bitmask[22];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10918_o = result_tmp[22];
  assign n10919_o = n10538_o[22];
  assign n10920_o = n10536_o[22];
  assign n10921_o = n10533_o[22];
  assign n10922_o = n10534_o[22];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10923_o = bf_bchg ? n10921_o : n10922_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10924_o = bf_ins ? n10920_o : n10923_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10925_o = bf_bset ? n10919_o : n10924_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10926_o = n10917_o ? n10918_o : n10925_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10934_o = shifted_bitmask[23];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10935_o = result_tmp[23];
  assign n10936_o = n10538_o[23];
  assign n10937_o = n10536_o[23];
  assign n10938_o = n10533_o[23];
  assign n10939_o = n10534_o[23];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10940_o = bf_bchg ? n10938_o : n10939_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10941_o = bf_ins ? n10937_o : n10940_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10942_o = bf_bset ? n10936_o : n10941_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10943_o = n10934_o ? n10935_o : n10942_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10951_o = shifted_bitmask[24];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10952_o = result_tmp[24];
  assign n10953_o = n10538_o[24];
  assign n10954_o = n10536_o[24];
  assign n10955_o = n10533_o[24];
  assign n10956_o = n10534_o[24];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10957_o = bf_bchg ? n10955_o : n10956_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10958_o = bf_ins ? n10954_o : n10957_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10959_o = bf_bset ? n10953_o : n10958_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10960_o = n10951_o ? n10952_o : n10959_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10968_o = shifted_bitmask[25];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10969_o = result_tmp[25];
  assign n10970_o = n10538_o[25];
  assign n10971_o = n10536_o[25];
  assign n10972_o = n10533_o[25];
  assign n10973_o = n10534_o[25];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10974_o = bf_bchg ? n10972_o : n10973_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10975_o = bf_ins ? n10971_o : n10974_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10976_o = bf_bset ? n10970_o : n10975_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10977_o = n10968_o ? n10969_o : n10976_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n10985_o = shifted_bitmask[26];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n10986_o = result_tmp[26];
  assign n10987_o = n10538_o[26];
  assign n10988_o = n10536_o[26];
  assign n10989_o = n10533_o[26];
  assign n10990_o = n10534_o[26];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n10991_o = bf_bchg ? n10989_o : n10990_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n10992_o = bf_ins ? n10988_o : n10991_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n10993_o = bf_bset ? n10987_o : n10992_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n10994_o = n10985_o ? n10986_o : n10993_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11002_o = shifted_bitmask[27];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11003_o = result_tmp[27];
  assign n11004_o = n10538_o[27];
  assign n11005_o = n10536_o[27];
  assign n11006_o = n10533_o[27];
  assign n11007_o = n10534_o[27];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11008_o = bf_bchg ? n11006_o : n11007_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11009_o = bf_ins ? n11005_o : n11008_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11010_o = bf_bset ? n11004_o : n11009_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11011_o = n11002_o ? n11003_o : n11010_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11019_o = shifted_bitmask[28];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11020_o = result_tmp[28];
  assign n11021_o = n10538_o[28];
  assign n11022_o = n10536_o[28];
  assign n11023_o = n10533_o[28];
  assign n11024_o = n10534_o[28];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11025_o = bf_bchg ? n11023_o : n11024_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11026_o = bf_ins ? n11022_o : n11025_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11027_o = bf_bset ? n11021_o : n11026_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11028_o = n11019_o ? n11020_o : n11027_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11036_o = shifted_bitmask[29];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11037_o = result_tmp[29];
  assign n11038_o = n10538_o[29];
  assign n11039_o = n10536_o[29];
  assign n11040_o = n10533_o[29];
  assign n11041_o = n10534_o[29];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11042_o = bf_bchg ? n11040_o : n11041_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11043_o = bf_ins ? n11039_o : n11042_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11044_o = bf_bset ? n11038_o : n11043_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11045_o = n11036_o ? n11037_o : n11044_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11053_o = shifted_bitmask[30];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11054_o = result_tmp[30];
  assign n11055_o = n10538_o[30];
  assign n11056_o = n10536_o[30];
  assign n11057_o = n10533_o[30];
  assign n11058_o = n10534_o[30];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11059_o = bf_bchg ? n11057_o : n11058_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11060_o = bf_ins ? n11056_o : n11059_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11061_o = bf_bset ? n11055_o : n11060_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11062_o = n11053_o ? n11054_o : n11061_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11070_o = shifted_bitmask[31];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11071_o = result_tmp[31];
  assign n11072_o = n10538_o[31];
  assign n11073_o = n10536_o[31];
  assign n11074_o = n10533_o[31];
  assign n11075_o = n10534_o[31];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11076_o = bf_bchg ? n11074_o : n11075_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11077_o = bf_ins ? n11073_o : n11076_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11078_o = bf_bset ? n11072_o : n11077_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11079_o = n11070_o ? n11071_o : n11078_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11087_o = shifted_bitmask[32];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11088_o = result_tmp[32];
  assign n11089_o = n10538_o[32];
  assign n11090_o = n10536_o[32];
  assign n11091_o = n10533_o[32];
  assign n11092_o = n10534_o[32];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11093_o = bf_bchg ? n11091_o : n11092_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11094_o = bf_ins ? n11090_o : n11093_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11095_o = bf_bset ? n11089_o : n11094_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11096_o = n11087_o ? n11088_o : n11095_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11104_o = shifted_bitmask[33];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11105_o = result_tmp[33];
  assign n11106_o = n10538_o[33];
  assign n11107_o = n10536_o[33];
  assign n11108_o = n10533_o[33];
  assign n11109_o = n10534_o[33];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11110_o = bf_bchg ? n11108_o : n11109_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11111_o = bf_ins ? n11107_o : n11110_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11112_o = bf_bset ? n11106_o : n11111_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11113_o = n11104_o ? n11105_o : n11112_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11121_o = shifted_bitmask[34];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11122_o = result_tmp[34];
  assign n11123_o = n10538_o[34];
  assign n11124_o = n10536_o[34];
  assign n11125_o = n10533_o[34];
  assign n11126_o = n10534_o[34];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11127_o = bf_bchg ? n11125_o : n11126_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11128_o = bf_ins ? n11124_o : n11127_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11129_o = bf_bset ? n11123_o : n11128_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11130_o = n11121_o ? n11122_o : n11129_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11138_o = shifted_bitmask[35];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11139_o = result_tmp[35];
  assign n11140_o = n10538_o[35];
  assign n11141_o = n10536_o[35];
  assign n11142_o = n10533_o[35];
  assign n11143_o = n10534_o[35];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11144_o = bf_bchg ? n11142_o : n11143_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11145_o = bf_ins ? n11141_o : n11144_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11146_o = bf_bset ? n11140_o : n11145_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11147_o = n11138_o ? n11139_o : n11146_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11155_o = shifted_bitmask[36];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11156_o = result_tmp[36];
  assign n11157_o = n10538_o[36];
  assign n11158_o = n10536_o[36];
  assign n11159_o = n10533_o[36];
  assign n11160_o = n10534_o[36];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11161_o = bf_bchg ? n11159_o : n11160_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11162_o = bf_ins ? n11158_o : n11161_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11163_o = bf_bset ? n11157_o : n11162_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11164_o = n11155_o ? n11156_o : n11163_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11172_o = shifted_bitmask[37];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11173_o = result_tmp[37];
  assign n11174_o = n10538_o[37];
  assign n11175_o = n10536_o[37];
  assign n11176_o = n10533_o[37];
  assign n11177_o = n10534_o[37];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11178_o = bf_bchg ? n11176_o : n11177_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11179_o = bf_ins ? n11175_o : n11178_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11180_o = bf_bset ? n11174_o : n11179_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11181_o = n11172_o ? n11173_o : n11180_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11189_o = shifted_bitmask[38];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11190_o = result_tmp[38];
  assign n11191_o = n10538_o[38];
  assign n11192_o = n10536_o[38];
  assign n11193_o = n10533_o[38];
  assign n11194_o = n10534_o[38];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11195_o = bf_bchg ? n11193_o : n11194_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11196_o = bf_ins ? n11192_o : n11195_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11197_o = bf_bset ? n11191_o : n11196_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11198_o = n11189_o ? n11190_o : n11197_o;
  assign n11199_o = n10538_o[39];
  assign n11200_o = n10536_o[39];
  assign n11201_o = n10533_o[39];
  assign n11202_o = n10534_o[39];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n11203_o = bf_bchg ? n11201_o : n11202_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n11204_o = bf_ins ? n11200_o : n11203_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n11205_o = bf_bset ? n11199_o : n11204_o;
  /* ../TG68K.C/TG68K_ALU.vhd:591:43  */
  assign n11206_o = shifted_bitmask[39];
  /* ../TG68K.C/TG68K_ALU.vhd:592:56  */
  assign n11207_o = result_tmp[39];
  /* ../TG68K.C/TG68K_ALU.vhd:591:25  */
  assign n11208_o = n11206_o ? n11207_o : n11205_o;
  /* ../TG68K.C/TG68K_ALU.vhd:598:36  */
  assign n11210_o = {1'b0, bitnr};
  /* ../TG68K.C/TG68K_ALU.vhd:598:43  */
  assign n11211_o = {5'b0, mask_not_zero};  //  uext
  /* ../TG68K.C/TG68K_ALU.vhd:598:43  */
  assign n11212_o = n11210_o + n11211_o;
  /* ../TG68K.C/TG68K_ALU.vhd:601:24  */
  assign n11213_o = mask[31:28];
  /* ../TG68K.C/TG68K_ALU.vhd:601:38  */
  assign n11215_o = n11213_o == 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:602:32  */
  assign n11216_o = mask[27:24];
  /* ../TG68K.C/TG68K_ALU.vhd:602:46  */
  assign n11218_o = n11216_o == 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:603:40  */
  assign n11219_o = mask[23:20];
  /* ../TG68K.C/TG68K_ALU.vhd:603:54  */
  assign n11221_o = n11219_o == 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:604:48  */
  assign n11222_o = mask[19:16];
  /* ../TG68K.C/TG68K_ALU.vhd:604:62  */
  assign n11224_o = n11222_o == 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:606:56  */
  assign n11226_o = mask[15:12];
  /* ../TG68K.C/TG68K_ALU.vhd:606:70  */
  assign n11228_o = n11226_o == 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:607:64  */
  assign n11229_o = mask[11:8];
  /* ../TG68K.C/TG68K_ALU.vhd:607:77  */
  assign n11231_o = n11229_o == 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:609:72  */
  assign n11233_o = mask[7:4];
  /* ../TG68K.C/TG68K_ALU.vhd:609:84  */
  assign n11235_o = n11233_o == 4'b0000;
  /* ../TG68K.C/TG68K_ALU.vhd:611:84  */
  assign n11237_o = mask[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:613:84  */
  assign n11238_o = mask[7:4];
  /* ../TG68K.C/TG68K_ALU.vhd:609:65  */
  assign n11239_o = n11235_o ? n11237_o : n11238_o;
  /* ../TG68K.C/TG68K_ALU.vhd:609:65  */
  assign n11241_o = n11235_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:616:76  */
  assign n11242_o = mask[11:8];
  /* ../TG68K.C/TG68K_ALU.vhd:607:57  */
  assign n11244_o = n11231_o ? n11239_o : n11242_o;
  assign n11245_o = {1'b0, n11241_o};
  assign n11246_o = n11245_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:607:57  */
  assign n11247_o = n11231_o ? n11246_o : 1'b0;
  assign n11248_o = n11245_o[1];
  /* ../TG68K.C/TG68K_ALU.vhd:607:57  */
  assign n11250_o = n11231_o ? n11248_o : 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:620:68  */
  assign n11251_o = mask[15:12];
  /* ../TG68K.C/TG68K_ALU.vhd:606:49  */
  assign n11252_o = n11228_o ? n11244_o : n11251_o;
  assign n11253_o = {n11250_o, n11247_o};
  /* ../TG68K.C/TG68K_ALU.vhd:606:49  */
  assign n11255_o = n11228_o ? n11253_o : 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:623:60  */
  assign n11256_o = mask[19:16];
  /* ../TG68K.C/TG68K_ALU.vhd:604:41  */
  assign n11259_o = n11224_o ? n11252_o : n11256_o;
  assign n11260_o = {1'b0, 1'b0};
  assign n11261_o = {1'b0, n11255_o};
  assign n11262_o = n11261_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:604:41  */
  assign n11263_o = n11224_o ? n11262_o : n11260_o;
  assign n11264_o = n11261_o[2];
  /* ../TG68K.C/TG68K_ALU.vhd:604:41  */
  assign n11266_o = n11224_o ? n11264_o : 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:628:52  */
  assign n11267_o = mask[23:20];
  /* ../TG68K.C/TG68K_ALU.vhd:603:33  */
  assign n11269_o = n11221_o ? n11259_o : n11267_o;
  assign n11270_o = {n11266_o, n11263_o};
  assign n11271_o = n11270_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:603:33  */
  assign n11273_o = n11221_o ? n11271_o : 1'b1;
  assign n11274_o = n11270_o[1];
  /* ../TG68K.C/TG68K_ALU.vhd:603:33  */
  assign n11275_o = n11221_o ? n11274_o : 1'b0;
  assign n11276_o = n11270_o[2];
  /* ../TG68K.C/TG68K_ALU.vhd:603:33  */
  assign n11278_o = n11221_o ? n11276_o : 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:632:44  */
  assign n11279_o = mask[27:24];
  /* ../TG68K.C/TG68K_ALU.vhd:602:25  */
  assign n11281_o = n11218_o ? n11269_o : n11279_o;
  assign n11282_o = {n11278_o, n11275_o, n11273_o};
  assign n11283_o = n11282_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:602:25  */
  assign n11284_o = n11218_o ? n11283_o : 1'b0;
  assign n11285_o = n11282_o[2:1];
  /* ../TG68K.C/TG68K_ALU.vhd:602:25  */
  assign n11287_o = n11218_o ? n11285_o : 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:636:36  */
  assign n11288_o = mask[31:28];
  /* ../TG68K.C/TG68K_ALU.vhd:601:17  */
  assign n11289_o = n11215_o ? n11281_o : n11288_o;
  assign n11290_o = {n11287_o, n11284_o};
  /* ../TG68K.C/TG68K_ALU.vhd:601:17  */
  assign n11292_o = n11215_o ? n11290_o : 3'b111;
  /* ../TG68K.C/TG68K_ALU.vhd:639:23  */
  assign n11295_o = mux[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:639:35  */
  assign n11297_o = n11295_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:641:31  */
  assign n11299_o = mux[1];
  /* ../TG68K.C/TG68K_ALU.vhd:641:34  */
  assign n11300_o = ~n11299_o;
  /* ../TG68K.C/TG68K_ALU.vhd:643:39  */
  assign n11302_o = mux[0];
  /* ../TG68K.C/TG68K_ALU.vhd:643:42  */
  assign n11303_o = ~n11302_o;
  /* ../TG68K.C/TG68K_ALU.vhd:643:33  */
  assign n11306_o = n11303_o ? 1'b0 : 1'b1;
  assign n11307_o = n11293_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:641:25  */
  assign n11308_o = n11300_o ? 1'b0 : n11307_o;
  /* ../TG68K.C/TG68K_ALU.vhd:641:25  */
  assign n11310_o = n11300_o ? n11306_o : 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:648:31  */
  assign n11311_o = mux[3];
  /* ../TG68K.C/TG68K_ALU.vhd:648:34  */
  assign n11312_o = ~n11311_o;
  assign n11314_o = n11293_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:648:25  */
  assign n11315_o = n11312_o ? 1'b0 : n11314_o;
  assign n11316_o = {1'b0, n11308_o};
  assign n11317_o = n11316_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:639:17  */
  assign n11318_o = n11297_o ? n11317_o : n11315_o;
  assign n11319_o = n11316_o[1];
  assign n11320_o = n11293_o[1];
  /* ../TG68K.C/TG68K_ALU.vhd:639:17  */
  assign n11321_o = n11297_o ? n11319_o : n11320_o;
  /* ../TG68K.C/TG68K_ALU.vhd:639:17  */
  assign n11324_o = n11297_o ? n11310_o : 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:659:32  */
  assign n11329_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:661:66  */
  assign n11330_o = op1out[7];
  /* ../TG68K.C/TG68K_ALU.vhd:660:25  */
  assign n11332_o = n11329_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:663:66  */
  assign n11333_o = op1out[15];
  /* ../TG68K.C/TG68K_ALU.vhd:662:25  */
  assign n11335_o = n11329_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:662:34  */
  assign n11337_o = n11329_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:662:34  */
  assign n11338_o = n11335_o | n11337_o;
  /* ../TG68K.C/TG68K_ALU.vhd:665:66  */
  assign n11339_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:664:25  */
  assign n11341_o = n11329_o == 2'b10;
  assign n11342_o = {n11341_o, n11338_o, n11332_o};
  /* ../TG68K.C/TG68K_ALU.vhd:659:17  */
  always @*
    case (n11342_o)
      3'b100: n11343_o = n11339_o;
      3'b010: n11343_o = n11333_o;
      3'b001: n11343_o = n11330_o;
      default: n11343_o = rot_rot;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:685:24  */
  assign n11361_o = exec[23];
  /* ../TG68K.C/TG68K_ALU.vhd:687:39  */
  assign n11362_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:688:36  */
  assign n11364_o = rot_bits == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:689:47  */
  assign n11365_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:688:25  */
  assign n11367_o = n11364_o ? n11365_o : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:694:38  */
  assign n11368_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:699:48  */
  assign n11371_o = op1out[0];
  /* ../TG68K.C/TG68K_ALU.vhd:700:48  */
  assign n11372_o = op1out[0];
  /* ../TG68K.C/TG68K_ALU.vhd:694:25  */
  assign n11392_o = n11368_o ? rot_rot : n11371_o;
  /* ../TG68K.C/TG68K_ALU.vhd:694:25  */
  assign n11393_o = n11368_o ? rot_rot : n11372_o;
  /* ../TG68K.C/TG68K_ALU.vhd:685:17  */
  assign n11396_o = n11361_o ? n11362_o : n11392_o;
  /* ../TG68K.C/TG68K_ALU.vhd:685:17  */
  assign n11397_o = n11361_o ? n11367_o : n11393_o;
  /* ../TG68K.C/TG68K_ALU.vhd:685:17  */
  assign n11398_o = n11361_o ? op1out : bsout;
  /* ../TG68K.C/TG68K_ALU.vhd:723:28  */
  assign n11403_o = rot_bits == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:724:40  */
  assign n11404_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:725:33  */
  assign n11406_o = n11404_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:727:33  */
  assign n11408_o = n11404_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:727:42  */
  assign n11410_o = n11404_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:727:42  */
  assign n11411_o = n11408_o | n11410_o;
  /* ../TG68K.C/TG68K_ALU.vhd:729:33  */
  assign n11413_o = n11404_o == 2'b10;
  assign n11414_o = {n11413_o, n11411_o, n11406_o};
  /* ../TG68K.C/TG68K_ALU.vhd:724:25  */
  always @*
    case (n11414_o)
      3'b100: n11419_o = 6'b100001;
      3'b010: n11419_o = 6'b010001;
      3'b001: n11419_o = 6'b001001;
      default: n11419_o = 6'b100000;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:734:40  */
  assign n11420_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:735:33  */
  assign n11422_o = n11420_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:737:33  */
  assign n11424_o = n11420_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:737:42  */
  assign n11426_o = n11420_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:737:42  */
  assign n11427_o = n11424_o | n11426_o;
  /* ../TG68K.C/TG68K_ALU.vhd:739:33  */
  assign n11429_o = n11420_o == 2'b10;
  assign n11430_o = {n11429_o, n11427_o, n11422_o};
  /* ../TG68K.C/TG68K_ALU.vhd:734:25  */
  always @*
    case (n11430_o)
      3'b100: n11435_o = 6'b100000;
      3'b010: n11435_o = 6'b010000;
      3'b001: n11435_o = 6'b001000;
      default: n11435_o = 6'b100000;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:723:17  */
  assign n11436_o = n11403_o ? n11419_o : n11435_o;
  /* ../TG68K.C/TG68K_ALU.vhd:745:30  */
  assign n11438_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:745:42  */
  assign n11440_o = n11438_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:745:55  */
  assign n11441_o = exec[81];
  /* ../TG68K.C/TG68K_ALU.vhd:745:64  */
  assign n11442_o = ~n11441_o;
  /* ../TG68K.C/TG68K_ALU.vhd:745:48  */
  assign n11443_o = n11440_o | n11442_o;
  /* ../TG68K.C/TG68K_ALU.vhd:747:33  */
  assign n11444_o = exe_opcode[5];
  /* ../TG68K.C/TG68K_ALU.vhd:748:43  */
  assign n11445_o = op2out[5:0];
  /* ../TG68K.C/TG68K_ALU.vhd:750:59  */
  assign n11446_o = exe_opcode[11:9];
  /* ../TG68K.C/TG68K_ALU.vhd:751:38  */
  assign n11447_o = exe_opcode[11:9];
  /* ../TG68K.C/TG68K_ALU.vhd:751:51  */
  assign n11449_o = n11447_o == 3'b000;
  /* ../TG68K.C/TG68K_ALU.vhd:751:25  */
  assign n11452_o = n11449_o ? 3'b001 : 3'b000;
  assign n11453_o = {n11452_o, n11446_o};
  /* ../TG68K.C/TG68K_ALU.vhd:747:17  */
  assign n11454_o = n11444_o ? n11445_o : n11453_o;
  /* ../TG68K.C/TG68K_ALU.vhd:745:17  */
  assign n11456_o = n11443_o ? 6'b000001 : n11454_o;
  /* ../TG68K.C/TG68K_ALU.vhd:762:29  */
  assign n11463_o = $unsigned(bs_shift) < $unsigned(ring);
  /* ../TG68K.C/TG68K_ALU.vhd:763:40  */
  assign n11464_o = ring - bs_shift;
  /* ../TG68K.C/TG68K_ALU.vhd:762:17  */
  assign n11466_o = n11463_o ? n11464_o : 6'b000000;
  /* ../TG68K.C/TG68K_ALU.vhd:765:45  */
  assign n11468_o = vector[30:0];
  /* ../TG68K.C/TG68K_ALU.vhd:765:38  */
  assign n11470_o = {1'b0, n11468_o};
  /* ../TG68K.C/TG68K_ALU.vhd:765:75  */
  assign n11471_o = vector[31:1];
  /* ../TG68K.C/TG68K_ALU.vhd:765:68  */
  assign n11473_o = {1'b0, n11471_o};
  /* ../TG68K.C/TG68K_ALU.vhd:765:60  */
  assign n11474_o = n11470_o ^ n11473_o;
  /* ../TG68K.C/TG68K_ALU.vhd:765:90  */
  assign n11475_o = {n11474_o, msb};
  /* ../TG68K.C/TG68K_ALU.vhd:766:32  */
  assign n11476_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:767:25  */
  assign n11479_o = n11476_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:769:25  */
  assign n11482_o = n11476_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:769:34  */
  assign n11484_o = n11476_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:769:34  */
  assign n11485_o = n11482_o | n11484_o;
  assign n11486_o = {n11485_o, n11479_o};
  assign n11487_o = n11475_o[8];
  /* ../TG68K.C/TG68K_ALU.vhd:766:17  */
  always @*
    case (n11486_o)
      2'b10: n11488_o = n11487_o;
      2'b01: n11488_o = 1'b0;
      default: n11488_o = n11487_o;
    endcase
  assign n11489_o = n11475_o[16];
  /* ../TG68K.C/TG68K_ALU.vhd:766:17  */
  always @*
    case (n11486_o)
      2'b10: n11490_o = 1'b0;
      2'b01: n11490_o = n11489_o;
      default: n11490_o = n11489_o;
    endcase
  assign n11492_o = n11475_o[7:0];
  assign n11493_o = n11475_o[32:17];
  assign n11494_o = n11475_o[15:9];
  /* ../TG68K.C/TG68K_ALU.vhd:773:56  */
  assign n11495_o = hot_msb[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:773:48  */
  assign n11497_o = {1'b0, n11495_o};
  /* ../TG68K.C/TG68K_ALU.vhd:773:42  */
  assign n11498_o = asl_over_xor - n11497_o;
  /* ../TG68K.C/TG68K_ALU.vhd:775:28  */
  assign n11500_o = rot_bits == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:775:48  */
  assign n11501_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:775:34  */
  assign n11502_o = n11500_o & n11501_o;
  /* ../TG68K.C/TG68K_ALU.vhd:776:45  */
  assign n11503_o = asl_over[32];
  /* ../TG68K.C/TG68K_ALU.vhd:776:33  */
  assign n11504_o = ~n11503_o;
  /* ../TG68K.C/TG68K_ALU.vhd:775:17  */
  assign n11506_o = n11502_o ? n11504_o : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:780:30  */
  assign n11508_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:780:33  */
  assign n11509_o = ~n11508_o;
  /* ../TG68K.C/TG68K_ALU.vhd:781:42  */
  assign n11510_o = result_bs[31];
  /* ../TG68K.C/TG68K_ALU.vhd:783:40  */
  assign n11511_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:785:58  */
  assign n11512_o = result_bs[8];
  /* ../TG68K.C/TG68K_ALU.vhd:784:33  */
  assign n11514_o = n11511_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:787:58  */
  assign n11515_o = result_bs[16];
  /* ../TG68K.C/TG68K_ALU.vhd:786:33  */
  assign n11517_o = n11511_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:786:42  */
  assign n11519_o = n11511_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:786:42  */
  assign n11520_o = n11517_o | n11519_o;
  /* ../TG68K.C/TG68K_ALU.vhd:789:58  */
  assign n11521_o = result_bs[32];
  /* ../TG68K.C/TG68K_ALU.vhd:788:33  */
  assign n11523_o = n11511_o == 2'b10;
  assign n11524_o = {n11523_o, n11520_o, n11514_o};
  /* ../TG68K.C/TG68K_ALU.vhd:783:25  */
  always @*
    case (n11524_o)
      3'b100: n11525_o = n11521_o;
      3'b010: n11525_o = n11515_o;
      3'b001: n11525_o = n11512_o;
      default: n11525_o = bs_c;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:780:17  */
  assign n11526_o = n11509_o ? n11510_o : n11525_o;
  /* ../TG68K.C/TG68K_ALU.vhd:795:28  */
  assign n11528_o = rot_bits == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:796:38  */
  assign n11529_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:797:40  */
  assign n11530_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:799:69  */
  assign n11531_o = result_bs[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:799:94  */
  assign n11532_o = result_bs[15:8];
  /* ../TG68K.C/TG68K_ALU.vhd:799:82  */
  assign n11533_o = n11531_o | n11532_o;
  /* ../TG68K.C/TG68K_ALU.vhd:800:52  */
  assign n11534_o = alu[7];
  /* ../TG68K.C/TG68K_ALU.vhd:798:33  */
  assign n11536_o = n11530_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:802:70  */
  assign n11537_o = result_bs[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:802:96  */
  assign n11538_o = result_bs[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:802:84  */
  assign n11539_o = n11537_o | n11538_o;
  /* ../TG68K.C/TG68K_ALU.vhd:803:52  */
  assign n11540_o = alu[15];
  /* ../TG68K.C/TG68K_ALU.vhd:801:33  */
  assign n11542_o = n11530_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:801:42  */
  assign n11544_o = n11530_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:801:42  */
  assign n11545_o = n11542_o | n11544_o;
  /* ../TG68K.C/TG68K_ALU.vhd:805:57  */
  assign n11546_o = result_bs[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:805:83  */
  assign n11547_o = result_bs[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:805:71  */
  assign n11548_o = n11546_o | n11547_o;
  /* ../TG68K.C/TG68K_ALU.vhd:806:52  */
  assign n11549_o = alu[31];
  /* ../TG68K.C/TG68K_ALU.vhd:804:33  */
  assign n11551_o = n11530_o == 2'b10;
  assign n11552_o = {n11551_o, n11545_o, n11536_o};
  assign n11553_o = n11539_o[7:0];
  assign n11554_o = n11548_o[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:797:25  */
  always @*
    case (n11552_o)
      3'b100: n11556_o = n11554_o;
      3'b010: n11556_o = n11553_o;
      3'b001: n11556_o = n11533_o;
      default: n11556_o = 8'bX;
    endcase
  assign n11557_o = n11539_o[15:8];
  assign n11558_o = n11548_o[15:8];
  /* ../TG68K.C/TG68K_ALU.vhd:797:25  */
  always @*
    case (n11552_o)
      3'b100: n11560_o = n11558_o;
      3'b010: n11560_o = n11557_o;
      3'b001: n11560_o = 8'bX;
      default: n11560_o = 8'bX;
    endcase
  assign n11561_o = n11548_o[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:797:25  */
  always @*
    case (n11552_o)
      3'b100: n11563_o = n11561_o;
      3'b010: n11563_o = 16'bX;
      3'b001: n11563_o = 16'bX;
      default: n11563_o = 16'bX;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:797:25  */
  always @*
    case (n11552_o)
      3'b100: n11564_o = n11549_o;
      3'b010: n11564_o = n11540_o;
      3'b001: n11564_o = n11534_o;
      default: n11564_o = n11526_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:809:38  */
  assign n11565_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:810:44  */
  assign n11566_o = alu[0];
  /* ../TG68K.C/TG68K_ALU.vhd:809:25  */
  assign n11567_o = n11565_o ? n11566_o : n11564_o;
  /* ../TG68K.C/TG68K_ALU.vhd:812:31  */
  assign n11569_o = rot_bits == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:813:40  */
  assign n11570_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:815:69  */
  assign n11571_o = result_bs[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:815:94  */
  assign n11572_o = result_bs[16:9];
  /* ../TG68K.C/TG68K_ALU.vhd:815:82  */
  assign n11573_o = n11571_o | n11572_o;
  /* ../TG68K.C/TG68K_ALU.vhd:816:58  */
  assign n11574_o = result_bs[8];
  /* ../TG68K.C/TG68K_ALU.vhd:816:74  */
  assign n11575_o = result_bs[17];
  /* ../TG68K.C/TG68K_ALU.vhd:816:62  */
  assign n11576_o = n11574_o | n11575_o;
  /* ../TG68K.C/TG68K_ALU.vhd:814:33  */
  assign n11578_o = n11570_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:818:70  */
  assign n11579_o = result_bs[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:818:96  */
  assign n11580_o = result_bs[32:17];
  /* ../TG68K.C/TG68K_ALU.vhd:818:84  */
  assign n11581_o = n11579_o | n11580_o;
  /* ../TG68K.C/TG68K_ALU.vhd:819:58  */
  assign n11582_o = result_bs[16];
  /* ../TG68K.C/TG68K_ALU.vhd:819:75  */
  assign n11583_o = result_bs[33];
  /* ../TG68K.C/TG68K_ALU.vhd:819:63  */
  assign n11584_o = n11582_o | n11583_o;
  /* ../TG68K.C/TG68K_ALU.vhd:817:33  */
  assign n11586_o = n11570_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:817:42  */
  assign n11588_o = n11570_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:817:42  */
  assign n11589_o = n11586_o | n11588_o;
  /* ../TG68K.C/TG68K_ALU.vhd:821:57  */
  assign n11590_o = result_bs[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:821:83  */
  assign n11591_o = result_bs[64:33];
  /* ../TG68K.C/TG68K_ALU.vhd:821:71  */
  assign n11592_o = n11590_o | n11591_o;
  /* ../TG68K.C/TG68K_ALU.vhd:822:58  */
  assign n11593_o = result_bs[32];
  /* ../TG68K.C/TG68K_ALU.vhd:822:75  */
  assign n11594_o = result_bs[65];
  /* ../TG68K.C/TG68K_ALU.vhd:822:63  */
  assign n11595_o = n11593_o | n11594_o;
  /* ../TG68K.C/TG68K_ALU.vhd:820:33  */
  assign n11597_o = n11570_o == 2'b10;
  assign n11598_o = {n11597_o, n11589_o, n11578_o};
  assign n11599_o = n11581_o[7:0];
  assign n11600_o = n11592_o[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:813:25  */
  always @*
    case (n11598_o)
      3'b100: n11602_o = n11600_o;
      3'b010: n11602_o = n11599_o;
      3'b001: n11602_o = n11573_o;
      default: n11602_o = 8'bX;
    endcase
  assign n11603_o = n11581_o[15:8];
  assign n11604_o = n11592_o[15:8];
  /* ../TG68K.C/TG68K_ALU.vhd:813:25  */
  always @*
    case (n11598_o)
      3'b100: n11606_o = n11604_o;
      3'b010: n11606_o = n11603_o;
      3'b001: n11606_o = 8'bX;
      default: n11606_o = 8'bX;
    endcase
  assign n11607_o = n11592_o[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:813:25  */
  always @*
    case (n11598_o)
      3'b100: n11609_o = n11607_o;
      3'b010: n11609_o = 16'bX;
      3'b001: n11609_o = 16'bX;
      default: n11609_o = 16'bX;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:813:25  */
  always @*
    case (n11598_o)
      3'b100: n11610_o = n11595_o;
      3'b010: n11610_o = n11584_o;
      3'b001: n11610_o = n11576_o;
      default: n11610_o = n11526_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:826:38  */
  assign n11611_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:826:41  */
  assign n11612_o = ~n11611_o;
  /* ../TG68K.C/TG68K_ALU.vhd:827:49  */
  assign n11613_o = result_bs[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:829:49  */
  assign n11614_o = result_bs[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:826:25  */
  assign n11615_o = n11612_o ? n11613_o : n11614_o;
  assign n11616_o = {n11609_o, n11606_o, n11602_o};
  /* ../TG68K.C/TG68K_ALU.vhd:812:17  */
  assign n11617_o = n11569_o ? n11616_o : n11615_o;
  /* ../TG68K.C/TG68K_ALU.vhd:812:17  */
  assign n11618_o = n11569_o ? n11610_o : n11526_o;
  assign n11619_o = {n11563_o, n11560_o, n11556_o};
  /* ../TG68K.C/TG68K_ALU.vhd:795:17  */
  assign n11620_o = n11528_o ? n11619_o : n11617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:795:17  */
  assign n11622_o = n11528_o ? n11567_o : n11618_o;
  /* ../TG68K.C/TG68K_ALU.vhd:795:17  */
  assign n11623_o = n11528_o ? n11529_o : bs_c;
  /* ../TG68K.C/TG68K_ALU.vhd:833:29  */
  assign n11625_o = bs_shift == 6'b000000;
  /* ../TG68K.C/TG68K_ALU.vhd:834:36  */
  assign n11627_o = rot_bits == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:835:46  */
  assign n11628_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:834:25  */
  assign n11630_o = n11627_o ? n11628_o : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:839:38  */
  assign n11631_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:833:17  */
  assign n11633_o = n11625_o ? 1'b0 : n11506_o;
  /* ../TG68K.C/TG68K_ALU.vhd:833:17  */
  assign n11634_o = n11625_o ? n11630_o : n11622_o;
  /* ../TG68K.C/TG68K_ALU.vhd:833:17  */
  assign n11635_o = n11625_o ? n11631_o : n11623_o;
  /* ../TG68K.C/TG68K_ALU.vhd:848:45  */
  assign n11637_o = bs_shift == 6'b111111;
  /* ../TG68K.C/TG68K_ALU.vhd:850:48  */
  assign n11639_o = $unsigned(bs_shift) > $unsigned(6'b110101);
  /* ../TG68K.C/TG68K_ALU.vhd:851:66  */
  assign n11641_o = bs_shift - 6'b110110;
  /* ../TG68K.C/TG68K_ALU.vhd:852:48  */
  assign n11643_o = $unsigned(bs_shift) > $unsigned(6'b101100);
  /* ../TG68K.C/TG68K_ALU.vhd:853:66  */
  assign n11645_o = bs_shift - 6'b101101;
  /* ../TG68K.C/TG68K_ALU.vhd:854:48  */
  assign n11647_o = $unsigned(bs_shift) > $unsigned(6'b100011);
  /* ../TG68K.C/TG68K_ALU.vhd:855:66  */
  assign n11649_o = bs_shift - 6'b100100;
  /* ../TG68K.C/TG68K_ALU.vhd:856:48  */
  assign n11651_o = $unsigned(bs_shift) > $unsigned(6'b011010);
  /* ../TG68K.C/TG68K_ALU.vhd:857:66  */
  assign n11653_o = bs_shift - 6'b011011;
  /* ../TG68K.C/TG68K_ALU.vhd:858:48  */
  assign n11655_o = $unsigned(bs_shift) > $unsigned(6'b010001);
  /* ../TG68K.C/TG68K_ALU.vhd:859:66  */
  assign n11657_o = bs_shift - 6'b010010;
  /* ../TG68K.C/TG68K_ALU.vhd:860:48  */
  assign n11659_o = $unsigned(bs_shift) > $unsigned(6'b001000);
  /* ../TG68K.C/TG68K_ALU.vhd:861:66  */
  assign n11661_o = bs_shift - 6'b001001;
  /* ../TG68K.C/TG68K_ALU.vhd:860:33  */
  assign n11662_o = n11659_o ? n11661_o : bs_shift;
  /* ../TG68K.C/TG68K_ALU.vhd:858:33  */
  assign n11663_o = n11655_o ? n11657_o : n11662_o;
  /* ../TG68K.C/TG68K_ALU.vhd:856:33  */
  assign n11664_o = n11651_o ? n11653_o : n11663_o;
  /* ../TG68K.C/TG68K_ALU.vhd:854:33  */
  assign n11665_o = n11647_o ? n11649_o : n11664_o;
  /* ../TG68K.C/TG68K_ALU.vhd:852:33  */
  assign n11666_o = n11643_o ? n11645_o : n11665_o;
  /* ../TG68K.C/TG68K_ALU.vhd:850:33  */
  assign n11667_o = n11639_o ? n11641_o : n11666_o;
  /* ../TG68K.C/TG68K_ALU.vhd:848:33  */
  assign n11669_o = n11637_o ? 6'b000000 : n11667_o;
  /* ../TG68K.C/TG68K_ALU.vhd:847:25  */
  assign n11671_o = ring == 6'b001001;
  /* ../TG68K.C/TG68K_ALU.vhd:866:45  */
  assign n11673_o = $unsigned(bs_shift) > $unsigned(6'b110010);
  /* ../TG68K.C/TG68K_ALU.vhd:867:66  */
  assign n11675_o = bs_shift - 6'b110011;
  /* ../TG68K.C/TG68K_ALU.vhd:868:48  */
  assign n11677_o = $unsigned(bs_shift) > $unsigned(6'b100001);
  /* ../TG68K.C/TG68K_ALU.vhd:869:66  */
  assign n11679_o = bs_shift - 6'b100010;
  /* ../TG68K.C/TG68K_ALU.vhd:870:48  */
  assign n11681_o = $unsigned(bs_shift) > $unsigned(6'b010000);
  /* ../TG68K.C/TG68K_ALU.vhd:871:66  */
  assign n11683_o = bs_shift - 6'b010001;
  /* ../TG68K.C/TG68K_ALU.vhd:870:33  */
  assign n11684_o = n11681_o ? n11683_o : bs_shift;
  /* ../TG68K.C/TG68K_ALU.vhd:868:33  */
  assign n11685_o = n11677_o ? n11679_o : n11684_o;
  /* ../TG68K.C/TG68K_ALU.vhd:866:33  */
  assign n11686_o = n11673_o ? n11675_o : n11685_o;
  /* ../TG68K.C/TG68K_ALU.vhd:865:25  */
  assign n11688_o = ring == 6'b010001;
  /* ../TG68K.C/TG68K_ALU.vhd:876:45  */
  assign n11690_o = $unsigned(bs_shift) > $unsigned(6'b100000);
  /* ../TG68K.C/TG68K_ALU.vhd:877:66  */
  assign n11692_o = bs_shift - 6'b100001;
  /* ../TG68K.C/TG68K_ALU.vhd:876:33  */
  assign n11693_o = n11690_o ? n11692_o : bs_shift;
  /* ../TG68K.C/TG68K_ALU.vhd:875:25  */
  assign n11695_o = ring == 6'b100001;
  /* ../TG68K.C/TG68K_ALU.vhd:881:74  */
  assign n11696_o = bs_shift[2:0];
  /* ../TG68K.C/TG68K_ALU.vhd:881:64  */
  assign n11698_o = {3'b000, n11696_o};
  /* ../TG68K.C/TG68K_ALU.vhd:881:25  */
  assign n11700_o = ring == 6'b001000;
  /* ../TG68K.C/TG68K_ALU.vhd:882:74  */
  assign n11701_o = bs_shift[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:882:64  */
  assign n11703_o = {2'b00, n11701_o};
  /* ../TG68K.C/TG68K_ALU.vhd:882:25  */
  assign n11705_o = ring == 6'b010000;
  /* ../TG68K.C/TG68K_ALU.vhd:883:74  */
  assign n11706_o = bs_shift[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:883:64  */
  assign n11708_o = {1'b0, n11706_o};
  /* ../TG68K.C/TG68K_ALU.vhd:883:25  */
  assign n11710_o = ring == 6'b100000;
  assign n11711_o = {n11710_o, n11705_o, n11700_o, n11695_o, n11688_o, n11671_o};
  /* ../TG68K.C/TG68K_ALU.vhd:846:17  */
  always @*
    case (n11711_o)
      6'b100000: n11713_o = n11708_o;
      6'b010000: n11713_o = n11703_o;
      6'b001000: n11713_o = n11698_o;
      6'b000100: n11713_o = n11693_o;
      6'b000010: n11713_o = n11686_o;
      6'b000001: n11713_o = n11669_o;
      default: n11713_o = 6'b000000;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:888:30  */
  assign n11714_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:888:33  */
  assign n11715_o = ~n11714_o;
  /* ../TG68K.C/TG68K_ALU.vhd:889:39  */
  assign n11716_o = ring - bs_shift_mod;
  /* ../TG68K.C/TG68K_ALU.vhd:888:17  */
  assign n11717_o = n11715_o ? n11716_o : bs_shift_mod;
  /* ../TG68K.C/TG68K_ALU.vhd:891:28  */
  assign n11718_o = rot_bits[1];
  /* ../TG68K.C/TG68K_ALU.vhd:891:31  */
  assign n11719_o = ~n11718_o;
  /* ../TG68K.C/TG68K_ALU.vhd:892:38  */
  assign n11720_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:892:41  */
  assign n11721_o = ~n11720_o;
  /* ../TG68K.C/TG68K_ALU.vhd:893:45  */
  assign n11723_o = 6'b100000 - bs_shift_mod;
  /* ../TG68K.C/TG68K_ALU.vhd:892:25  */
  assign n11724_o = n11721_o ? n11723_o : n11717_o;
  /* ../TG68K.C/TG68K_ALU.vhd:895:37  */
  assign n11725_o = bs_shift == ring;
  /* ../TG68K.C/TG68K_ALU.vhd:896:46  */
  assign n11726_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:896:49  */
  assign n11727_o = ~n11726_o;
  /* ../TG68K.C/TG68K_ALU.vhd:897:53  */
  assign n11729_o = 6'b100000 - ring;
  /* ../TG68K.C/TG68K_ALU.vhd:896:33  */
  assign n11730_o = n11727_o ? n11729_o : ring;
  /* ../TG68K.C/TG68K_ALU.vhd:895:25  */
  assign n11731_o = n11725_o ? n11730_o : n11724_o;
  /* ../TG68K.C/TG68K_ALU.vhd:902:37  */
  assign n11732_o = $unsigned(bs_shift) > $unsigned(ring);
  /* ../TG68K.C/TG68K_ALU.vhd:903:46  */
  assign n11733_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:903:49  */
  assign n11734_o = ~n11733_o;
  /* ../TG68K.C/TG68K_ALU.vhd:907:55  */
  assign n11736_o = ring + 6'b000001;
  /* ../TG68K.C/TG68K_ALU.vhd:903:33  */
  assign n11738_o = n11734_o ? 6'b000000 : n11736_o;
  /* ../TG68K.C/TG68K_ALU.vhd:891:17  */
  assign n11740_o = n11744_o ? 1'b0 : n11634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:902:25  */
  assign n11741_o = n11732_o ? n11738_o : n11731_o;
  /* ../TG68K.C/TG68K_ALU.vhd:902:25  */
  assign n11742_o = n11732_o & n11734_o;
  /* ../TG68K.C/TG68K_ALU.vhd:891:17  */
  assign n11743_o = n11719_o ? n11741_o : n11717_o;
  /* ../TG68K.C/TG68K_ALU.vhd:891:17  */
  assign n11744_o = n11719_o & n11742_o;
  /* ../TG68K.C/TG68K_ALU.vhd:915:50  */
  assign n11745_o = asr_sign[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:915:74  */
  assign n11746_o = hot_msb[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:915:64  */
  assign n11747_o = n11745_o | n11746_o;
  assign n11749_o = n11748_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:916:28  */
  assign n11751_o = rot_bits == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:916:48  */
  assign n11752_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:916:51  */
  assign n11753_o = ~n11752_o;
  /* ../TG68K.C/TG68K_ALU.vhd:916:34  */
  assign n11754_o = n11751_o & n11753_o;
  /* ../TG68K.C/TG68K_ALU.vhd:916:56  */
  assign n11755_o = n11754_o & msb;
  /* ../TG68K.C/TG68K_ALU.vhd:917:49  */
  assign n11756_o = asr_sign[32:1];
  /* ../TG68K.C/TG68K_ALU.vhd:917:38  */
  assign n11757_o = alu | n11756_o;
  /* ../TG68K.C/TG68K_ALU.vhd:918:37  */
  assign n11758_o = $unsigned(bs_shift) > $unsigned(ring);
  /* ../TG68K.C/TG68K_ALU.vhd:916:17  */
  assign n11760_o = n11762_o ? 1'b1 : n11740_o;
  /* ../TG68K.C/TG68K_ALU.vhd:916:17  */
  assign n11762_o = n11755_o & n11758_o;
  /* ../TG68K.C/TG68K_ALU.vhd:923:43  */
  assign n11764_o = {1'b0, op1out};
  /* ../TG68K.C/TG68K_ALU.vhd:924:32  */
  assign n11765_o = exe_opcode[7:6];
  /* ../TG68K.C/TG68K_ALU.vhd:926:46  */
  assign n11766_o = op1out[7];
  /* ../TG68K.C/TG68K_ALU.vhd:929:44  */
  assign n11770_o = rot_bits == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:930:59  */
  assign n11771_o = n12543_q[4];
  assign n11772_o = n11767_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:929:33  */
  assign n11773_o = n11770_o ? n11771_o : n11772_o;
  assign n11774_o = n11767_o[23:1];
  /* ../TG68K.C/TG68K_ALU.vhd:925:25  */
  assign n11776_o = n11765_o == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:933:46  */
  assign n11777_o = op1out[15];
  /* ../TG68K.C/TG68K_ALU.vhd:936:44  */
  assign n11781_o = rot_bits == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:937:60  */
  assign n11782_o = n12543_q[4];
  assign n11783_o = n11778_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:936:33  */
  assign n11784_o = n11781_o ? n11782_o : n11783_o;
  assign n11785_o = n11778_o[15:1];
  /* ../TG68K.C/TG68K_ALU.vhd:932:25  */
  assign n11787_o = n11765_o == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:932:34  */
  assign n11789_o = n11765_o == 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:932:34  */
  assign n11790_o = n11787_o | n11789_o;
  /* ../TG68K.C/TG68K_ALU.vhd:940:46  */
  assign n11791_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:941:44  */
  assign n11793_o = rot_bits == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:942:60  */
  assign n11794_o = n12543_q[4];
  assign n11795_o = n11764_o[32];
  /* ../TG68K.C/TG68K_ALU.vhd:941:33  */
  assign n11796_o = n11793_o ? n11794_o : n11795_o;
  /* ../TG68K.C/TG68K_ALU.vhd:939:25  */
  assign n11798_o = n11765_o == 2'b10;
  assign n11799_o = {n11798_o, n11790_o, n11776_o};
  assign n11800_o = n11764_o[8];
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11801_o = n11800_o;
      3'b010: n11801_o = n11800_o;
      3'b001: n11801_o = n11773_o;
      default: n11801_o = n11800_o;
    endcase
  assign n11802_o = n11774_o[6:0];
  assign n11803_o = n11764_o[15:9];
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11804_o = n11803_o;
      3'b010: n11804_o = n11803_o;
      3'b001: n11804_o = n11802_o;
      default: n11804_o = n11803_o;
    endcase
  assign n11805_o = n11774_o[7];
  assign n11806_o = n11764_o[16];
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11807_o = n11806_o;
      3'b010: n11807_o = n11784_o;
      3'b001: n11807_o = n11805_o;
      default: n11807_o = n11806_o;
    endcase
  assign n11808_o = n11774_o[22:8];
  assign n11809_o = n11764_o[31:17];
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11810_o = n11809_o;
      3'b010: n11810_o = n11785_o;
      3'b001: n11810_o = n11808_o;
      default: n11810_o = n11809_o;
    endcase
  assign n11811_o = n11764_o[32];
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11812_o = n11796_o;
      3'b010: n11812_o = n11811_o;
      3'b001: n11812_o = n11811_o;
      default: n11812_o = n11811_o;
    endcase
  assign n11814_o = n11764_o[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11818_o = n11791_o;
      3'b010: n11818_o = n11777_o;
      3'b001: n11818_o = n11766_o;
      default: n11818_o = msb;
    endcase
  assign n11819_o = n11768_o[7:0];
  assign n11820_o = n11757_o[15:8];
  assign n11821_o = alu[15:8];
  /* ../TG68K.C/TG68K_ALU.vhd:916:17  */
  assign n11822_o = n11755_o ? n11820_o : n11821_o;
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11823_o = n11822_o;
      3'b010: n11823_o = n11822_o;
      3'b001: n11823_o = n11819_o;
      default: n11823_o = n11822_o;
    endcase
  assign n11824_o = n11768_o[23:8];
  assign n11825_o = n11757_o[31:16];
  assign n11826_o = alu[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:916:17  */
  assign n11827_o = n11755_o ? n11825_o : n11826_o;
  /* ../TG68K.C/TG68K_ALU.vhd:924:17  */
  always @*
    case (n11799_o)
      3'b100: n11828_o = n11827_o;
      3'b010: n11828_o = 16'b0000000000000000;
      3'b001: n11828_o = n11824_o;
      default: n11828_o = n11827_o;
    endcase
  assign n11832_o = n11757_o[7:0];
  assign n11833_o = alu[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:916:17  */
  assign n11834_o = n11755_o ? n11832_o : n11833_o;
  /* ../TG68K.C/TG68K_ALU.vhd:946:71  */
  assign n11836_o = {33'b000000000000000000000000000000000, vector};
  /* ../TG68K.C/TG68K_ALU.vhd:946:84  */
  assign n11837_o = {25'b0, bit_nr};  //  uext
  /* ../TG68K.C/TG68K_ALU.vhd:946:80  */
  assign n11838_o = {1'b0, n11837_o};  //  uext
  /* ../TG68K.C/TG68K_ALU.vhd:946:80  */
  assign n11839_o = n11836_o << n11838_o;
  /* ../TG68K.C/TG68K_ALU.vhd:957:24  */
  assign n11843_o = exec[17];
  /* ../TG68K.C/TG68K_ALU.vhd:958:58  */
  assign n11844_o = last_data_read[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:958:40  */
  assign n11845_o = n12543_q & n11844_o;
  /* ../TG68K.C/TG68K_ALU.vhd:959:27  */
  assign n11846_o = exec[18];
  /* ../TG68K.C/TG68K_ALU.vhd:960:58  */
  assign n11847_o = last_data_read[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:960:40  */
  assign n11848_o = n12543_q ^ n11847_o;
  /* ../TG68K.C/TG68K_ALU.vhd:961:27  */
  assign n11849_o = exec[19];
  /* ../TG68K.C/TG68K_ALU.vhd:962:57  */
  assign n11850_o = last_data_read[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:962:40  */
  assign n11851_o = n12543_q | n11850_o;
  /* ../TG68K.C/TG68K_ALU.vhd:964:40  */
  assign n11852_o = op2out[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:961:17  */
  assign n11853_o = n11849_o ? n11851_o : n11852_o;
  /* ../TG68K.C/TG68K_ALU.vhd:959:17  */
  assign n11854_o = n11846_o ? n11848_o : n11853_o;
  /* ../TG68K.C/TG68K_ALU.vhd:957:17  */
  assign n11855_o = n11843_o ? n11845_o : n11854_o;
  /* ../TG68K.C/TG68K_ALU.vhd:971:24  */
  assign n11856_o = exec[28];
  /* ../TG68K.C/TG68K_ALU.vhd:971:50  */
  assign n11857_o = n12543_q[2];
  /* ../TG68K.C/TG68K_ALU.vhd:971:53  */
  assign n11858_o = ~n11857_o;
  /* ../TG68K.C/TG68K_ALU.vhd:971:41  */
  assign n11859_o = n11856_o & n11858_o;
  /* ../TG68K.C/TG68K_ALU.vhd:973:28  */
  assign n11860_o = op1in[7:0];
  /* ../TG68K.C/TG68K_ALU.vhd:973:40  */
  assign n11862_o = n11860_o == 8'b00000000;
  /* ../TG68K.C/TG68K_ALU.vhd:975:33  */
  assign n11864_o = op1in[15:8];
  /* ../TG68K.C/TG68K_ALU.vhd:975:46  */
  assign n11866_o = n11864_o == 8'b00000000;
  /* ../TG68K.C/TG68K_ALU.vhd:977:41  */
  assign n11868_o = op1in[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:977:55  */
  assign n11870_o = n11868_o == 16'b0000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:977:33  */
  assign n11873_o = n11870_o ? 1'b1 : 1'b0;
  assign n11874_o = {n11873_o, 1'b1};
  /* ../TG68K.C/TG68K_ALU.vhd:975:25  */
  assign n11876_o = n11866_o ? n11874_o : 2'b00;
  assign n11877_o = {n11876_o, 1'b1};
  /* ../TG68K.C/TG68K_ALU.vhd:973:17  */
  assign n11879_o = n11862_o ? n11877_o : 3'b000;
  /* ../TG68K.C/TG68K_ALU.vhd:971:17  */
  assign n11881_o = n11859_o ? 3'b000 : n11879_o;
  /* ../TG68K.C/TG68K_ALU.vhd:984:32  */
  assign n11884_o = exe_datatype == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:985:43  */
  assign n11885_o = op1in[7];
  /* ../TG68K.C/TG68K_ALU.vhd:985:53  */
  assign n11886_o = flag_z[0];
  /* ../TG68K.C/TG68K_ALU.vhd:985:46  */
  assign n11887_o = {n11885_o, n11886_o};
  /* ../TG68K.C/TG68K_ALU.vhd:985:67  */
  assign n11888_o = addsub_ofl[0];
  /* ../TG68K.C/TG68K_ALU.vhd:985:56  */
  assign n11889_o = {n11887_o, n11888_o};
  /* ../TG68K.C/TG68K_ALU.vhd:985:76  */
  assign n11890_o = n9786_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:985:70  */
  assign n11891_o = {n11889_o, n11890_o};
  /* ../TG68K.C/TG68K_ALU.vhd:986:32  */
  assign n11892_o = exec[12];
  /* ../TG68K.C/TG68K_ALU.vhd:986:53  */
  assign n11893_o = exec[13];
  /* ../TG68K.C/TG68K_ALU.vhd:986:46  */
  assign n11894_o = n11892_o | n11893_o;
  assign n11895_o = {vflag_a, bcd_a_carry};
  assign n11896_o = n11891_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:986:25  */
  assign n11897_o = n11894_o ? n11895_o : n11896_o;
  assign n11898_o = n11891_o[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:990:35  */
  assign n11900_o = exe_datatype == 2'b10;
  /* ../TG68K.C/TG68K_ALU.vhd:990:48  */
  assign n11901_o = exec[10];
  /* ../TG68K.C/TG68K_ALU.vhd:990:41  */
  assign n11902_o = n11900_o | n11901_o;
  /* ../TG68K.C/TG68K_ALU.vhd:991:43  */
  assign n11903_o = op1in[31];
  /* ../TG68K.C/TG68K_ALU.vhd:991:54  */
  assign n11904_o = flag_z[2];
  /* ../TG68K.C/TG68K_ALU.vhd:991:47  */
  assign n11905_o = {n11903_o, n11904_o};
  /* ../TG68K.C/TG68K_ALU.vhd:991:68  */
  assign n11906_o = addsub_ofl[2];
  /* ../TG68K.C/TG68K_ALU.vhd:991:57  */
  assign n11907_o = {n11905_o, n11906_o};
  /* ../TG68K.C/TG68K_ALU.vhd:991:77  */
  assign n11908_o = n9786_o[2];
  /* ../TG68K.C/TG68K_ALU.vhd:991:71  */
  assign n11909_o = {n11907_o, n11908_o};
  /* ../TG68K.C/TG68K_ALU.vhd:993:43  */
  assign n11910_o = op1in[15];
  /* ../TG68K.C/TG68K_ALU.vhd:993:54  */
  assign n11911_o = flag_z[1];
  /* ../TG68K.C/TG68K_ALU.vhd:993:47  */
  assign n11912_o = {n11910_o, n11911_o};
  /* ../TG68K.C/TG68K_ALU.vhd:993:68  */
  assign n11913_o = addsub_ofl[1];
  /* ../TG68K.C/TG68K_ALU.vhd:993:57  */
  assign n11914_o = {n11912_o, n11913_o};
  /* ../TG68K.C/TG68K_ALU.vhd:993:77  */
  assign n11915_o = n9786_o[1];
  /* ../TG68K.C/TG68K_ALU.vhd:993:71  */
  assign n11916_o = {n11914_o, n11915_o};
  /* ../TG68K.C/TG68K_ALU.vhd:990:17  */
  assign n11917_o = n11902_o ? n11909_o : n11916_o;
  assign n11918_o = {n11898_o, n11897_o};
  /* ../TG68K.C/TG68K_ALU.vhd:984:17  */
  assign n11919_o = n11884_o ? n11918_o : n11917_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1000:40  */
  assign n11921_o = exec[59];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:55  */
  assign n11922_o = n11921_o | set_stop;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:40  */
  assign n11925_o = exec[60];
  /* ../TG68K.C/TG68K_ALU.vhd:1007:40  */
  assign n11928_o = exec[9];
  /* ../TG68K.C/TG68K_ALU.vhd:1007:66  */
  assign n11929_o = ~decodeopc;
  /* ../TG68K.C/TG68K_ALU.vhd:1007:53  */
  assign n11930_o = n11928_o & n11929_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1008:65  */
  assign n11931_o = set_flags[3];
  /* ../TG68K.C/TG68K_ALU.vhd:1008:69  */
  assign n11932_o = n11931_o ^ rot_rot;
  /* ../TG68K.C/TG68K_ALU.vhd:1008:82  */
  assign n11933_o = n11932_o | asl_vflag;
  /* ../TG68K.C/TG68K_ALU.vhd:1007:33  */
  assign n11935_o = n11930_o ? n11933_o : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:1012:40  */
  assign n11936_o = exec[51];
  /* ../TG68K.C/TG68K_ALU.vhd:1015:56  */
  assign n11938_o = micro_state == 7'b0110011;
  /* ../TG68K.C/TG68K_ALU.vhd:1017:62  */
  assign n11939_o = exe_opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:1017:65  */
  assign n11940_o = ~n11939_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1019:92  */
  assign n11941_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1019:82  */
  assign n11942_o = ~n11941_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1019:81  */
  assign n11944_o = {1'b0, n11942_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1019:96  */
  assign n11946_o = {n11944_o, 2'b00};
  /* ../TG68K.C/TG68K_ALU.vhd:1017:49  */
  assign n11948_o = n11940_o ? n11946_o : 4'b0100;
  assign n11949_o = data_read[3:0];
  assign n11950_o = data_read[3:0];
  assign n11951_o = n12543_q[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n11952_o = n11922_o ? n11950_o : n11951_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n11953_o = n11925_o ? n11949_o : n11952_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1015:41  */
  assign n11954_o = n11938_o ? n11948_o : n11953_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1024:43  */
  assign n11955_o = exec[49];
  /* ../TG68K.C/TG68K_ALU.vhd:1024:53  */
  assign n11956_o = ~n11955_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1025:61  */
  assign n11957_o = n12543_q[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1026:48  */
  assign n11958_o = exec[3];
  /* ../TG68K.C/TG68K_ALU.vhd:1027:70  */
  assign n11959_o = set_flags[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1028:51  */
  assign n11960_o = exec[9];
  /* ../TG68K.C/TG68K_ALU.vhd:1028:76  */
  assign n11962_o = rot_bits != 2'b11;
  /* ../TG68K.C/TG68K_ALU.vhd:1028:64  */
  assign n11963_o = n11960_o & n11962_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1028:91  */
  assign n11964_o = exec[23];
  /* ../TG68K.C/TG68K_ALU.vhd:1028:100  */
  assign n11965_o = ~n11964_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1028:83  */
  assign n11966_o = n11963_o & n11965_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1030:51  */
  assign n11967_o = exec[81];
  assign n11968_o = data_read[4];
  assign n11969_o = data_read[4];
  assign n11970_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n11971_o = n11922_o ? n11969_o : n11970_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n11972_o = n11925_o ? n11968_o : n11971_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1030:41  */
  assign n11973_o = n11967_o ? bs_x : n11972_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1028:41  */
  assign n11974_o = n11966_o ? rot_x : n11973_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1026:41  */
  assign n11975_o = n11958_o ? n11959_o : n11974_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1034:49  */
  assign n11976_o = exec[8];
  /* ../TG68K.C/TG68K_ALU.vhd:1034:65  */
  assign n11977_o = exec[86];
  /* ../TG68K.C/TG68K_ALU.vhd:1034:58  */
  assign n11978_o = n11976_o | n11977_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1036:51  */
  assign n11979_o = exec[21];
  /* ../TG68K.C/TG68K_ALU.vhd:1036:65  */
  assign n11981_o = n11979_o & 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:1039:65  */
  assign n11983_o = exe_opcode[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1039:74  */
  assign n11985_o = n11983_o | 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:1040:83  */
  assign n11986_o = op1in[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1040:94  */
  assign n11987_o = flag_z[1];
  /* ../TG68K.C/TG68K_ALU.vhd:1040:87  */
  assign n11988_o = {n11986_o, n11987_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1040:97  */
  assign n11990_o = {n11988_o, 2'b00};
  /* ../TG68K.C/TG68K_ALU.vhd:1042:83  */
  assign n11991_o = op1in[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1042:94  */
  assign n11992_o = flag_z[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1042:87  */
  assign n11993_o = {n11991_o, n11992_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1042:97  */
  assign n11995_o = {n11993_o, 2'b00};
  /* ../TG68K.C/TG68K_ALU.vhd:1039:49  */
  assign n11996_o = n11985_o ? n11990_o : n11995_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1037:49  */
  assign n11997_o = v_flag ? 4'b1010 : n11996_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1044:51  */
  assign n11998_o = exec[68];
  /* ../TG68K.C/TG68K_ALU.vhd:1044:72  */
  assign n12000_o = n11998_o & 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:1045:70  */
  assign n12001_o = set_flags[3];
  /* ../TG68K.C/TG68K_ALU.vhd:1046:70  */
  assign n12002_o = set_flags[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1046:83  */
  assign n12003_o = n12543_q[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1046:74  */
  assign n12004_o = n12002_o & n12003_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1049:51  */
  assign n12007_o = exec[67];
  /* ../TG68K.C/TG68K_ALU.vhd:1049:71  */
  assign n12009_o = n12007_o & 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:1050:70  */
  assign n12010_o = set_flags[3];
  /* ../TG68K.C/TG68K_ALU.vhd:1051:70  */
  assign n12011_o = set_flags[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:51  */
  assign n12013_o = exec[5];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:70  */
  assign n12014_o = exec[6];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:63  */
  assign n12015_o = n12013_o | n12014_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1054:90  */
  assign n12016_o = exec[7];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:83  */
  assign n12017_o = n12015_o | n12016_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1054:110  */
  assign n12018_o = exec[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:103  */
  assign n12019_o = n12017_o | n12018_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1054:131  */
  assign n12020_o = exec[1];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:124  */
  assign n12021_o = n12019_o | n12020_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1054:153  */
  assign n12022_o = exec[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:146  */
  assign n12023_o = n12021_o | n12022_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1054:174  */
  assign n12024_o = exec[75];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:167  */
  assign n12025_o = n12023_o | n12024_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1054:194  */
  assign n12026_o = exec[20];
  /* ../TG68K.C/TG68K_ALU.vhd:1054:208  */
  assign n12028_o = n12026_o & 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:1054:186  */
  assign n12029_o = n12025_o | n12028_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1057:56  */
  assign n12032_o = exec[75];
  assign n12033_o = set_flags[3];
  /* ../TG68K.C/TG68K_ALU.vhd:1057:49  */
  assign n12034_o = n12032_o ? bf_nflag : n12033_o;
  assign n12035_o = set_flags[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1060:51  */
  assign n12036_o = exec[9];
  /* ../TG68K.C/TG68K_ALU.vhd:1061:79  */
  assign n12037_o = set_flags[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:1063:60  */
  assign n12039_o = rot_bits == 2'b00;
  /* ../TG68K.C/TG68K_ALU.vhd:1063:81  */
  assign n12040_o = set_flags[3];
  /* ../TG68K.C/TG68K_ALU.vhd:1063:85  */
  assign n12041_o = n12040_o ^ rot_rot;
  /* ../TG68K.C/TG68K_ALU.vhd:1063:98  */
  assign n12042_o = n12041_o | asl_vflag;
  /* ../TG68K.C/TG68K_ALU.vhd:1063:66  */
  assign n12043_o = n12039_o & n12042_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1063:49  */
  assign n12046_o = n12043_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:1068:51  */
  assign n12047_o = exec[81];
  /* ../TG68K.C/TG68K_ALU.vhd:1069:79  */
  assign n12048_o = set_flags[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:1072:51  */
  assign n12049_o = exec[14];
  /* ../TG68K.C/TG68K_ALU.vhd:1073:61  */
  assign n12050_o = ~one_bit_in;
  /* ../TG68K.C/TG68K_ALU.vhd:1074:51  */
  assign n12051_o = exec[87];
  /* ../TG68K.C/TG68K_ALU.vhd:1079:63  */
  assign n12052_o = last_flags1[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1079:66  */
  assign n12053_o = ~n12052_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1080:74  */
  assign n12054_o = n12543_q[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1080:95  */
  assign n12055_o = set_flags[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1080:82  */
  assign n12056_o = ~n12055_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1080:116  */
  assign n12057_o = set_flags[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1080:103  */
  assign n12058_o = ~n12057_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1080:99  */
  assign n12059_o = n12056_o & n12058_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1080:78  */
  assign n12060_o = n12054_o | n12059_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1082:75  */
  assign n12061_o = n12543_q[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1082:92  */
  assign n12062_o = set_flags[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1082:79  */
  assign n12063_o = n12061_o ^ n12062_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1082:111  */
  assign n12064_o = n12543_q[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1082:102  */
  assign n12065_o = ~n12064_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1082:97  */
  assign n12066_o = n12063_o & n12065_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1082:132  */
  assign n12067_o = set_flags[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1082:119  */
  assign n12068_o = ~n12067_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1082:115  */
  assign n12069_o = n12066_o & n12068_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1079:49  */
  assign n12070_o = n12053_o ? n12060_o : n12069_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1085:66  */
  assign n12072_o = n12543_q[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1085:82  */
  assign n12073_o = set_flags[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1085:70  */
  assign n12074_o = n12072_o | n12073_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1086:76  */
  assign n12075_o = last_flags1[0];
  /* ../TG68K.C/TG68K_ALU.vhd:1086:61  */
  assign n12076_o = ~n12075_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1087:51  */
  assign n12077_o = exec[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1088:64  */
  assign n12079_o = exe_datatype == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:1089:75  */
  assign n12080_o = op1out[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1091:75  */
  assign n12081_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1088:49  */
  assign n12082_o = n12079_o ? n12080_o : n12081_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1093:58  */
  assign n12083_o = op1out[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1093:71  */
  assign n12085_o = n12083_o == 16'b0000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:1093:97  */
  assign n12087_o = exe_datatype == 2'b01;
  /* ../TG68K.C/TG68K_ALU.vhd:1093:112  */
  assign n12088_o = op1out[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1093:126  */
  assign n12090_o = n12088_o == 16'b0000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:1093:103  */
  assign n12091_o = n12087_o | n12090_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1093:80  */
  assign n12092_o = n12085_o & n12091_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1093:49  */
  assign n12095_o = n12092_o ? 1'b1 : 1'b0;
  assign n12098_o = {n12082_o, n12095_o, 1'b0, 1'b0};
  assign n12099_o = data_read[3:0];
  assign n12100_o = data_read[3:0];
  assign n12101_o = n12543_q[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n12102_o = n11922_o ? n12100_o : n12101_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n12103_o = n11925_o ? n12099_o : n12102_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1087:41  */
  assign n12104_o = n12077_o ? n12098_o : n12103_o;
  assign n12105_o = {n12076_o, n12074_o, 1'b0, n12070_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1074:41  */
  assign n12106_o = n12051_o ? n12105_o : n12104_o;
  assign n12107_o = n12106_o[1:0];
  assign n12108_o = data_read[1:0];
  assign n12109_o = data_read[1:0];
  assign n12110_o = n12543_q[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n12111_o = n11922_o ? n12109_o : n12110_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n12112_o = n11925_o ? n12108_o : n12111_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1072:41  */
  assign n12113_o = n12049_o ? n12112_o : n12107_o;
  assign n12114_o = n12106_o[2];
  /* ../TG68K.C/TG68K_ALU.vhd:1072:41  */
  assign n12115_o = n12049_o ? n12050_o : n12114_o;
  assign n12116_o = n12106_o[3];
  assign n12117_o = data_read[3];
  assign n12118_o = data_read[3];
  assign n12119_o = n12543_q[3];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n12120_o = n11922_o ? n12118_o : n12119_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n12121_o = n11925_o ? n12117_o : n12120_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1072:41  */
  assign n12122_o = n12049_o ? n12121_o : n12116_o;
  assign n12123_o = {n12122_o, n12115_o, n12113_o};
  assign n12124_o = {n12048_o, bs_v, bs_c};
  /* ../TG68K.C/TG68K_ALU.vhd:1068:41  */
  assign n12125_o = n12047_o ? n12124_o : n12123_o;
  assign n12126_o = {n12037_o, n12046_o, rot_c};
  /* ../TG68K.C/TG68K_ALU.vhd:1060:41  */
  assign n12127_o = n12036_o ? n12126_o : n12125_o;
  assign n12128_o = {n12034_o, n12035_o, 2'b00};
  /* ../TG68K.C/TG68K_ALU.vhd:1054:41  */
  assign n12129_o = n12029_o ? n12128_o : n12127_o;
  assign n12130_o = {n12010_o, n12011_o, set_mv_flag, 1'b0};
  /* ../TG68K.C/TG68K_ALU.vhd:1049:41  */
  assign n12131_o = n12009_o ? n12130_o : n12129_o;
  assign n12132_o = {n12001_o, n12004_o, 1'b0, 1'b0};
  /* ../TG68K.C/TG68K_ALU.vhd:1044:41  */
  assign n12133_o = n12000_o ? n12132_o : n12131_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1036:41  */
  assign n12134_o = n11981_o ? n11997_o : n12133_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1034:41  */
  assign n12135_o = n11978_o ? set_flags : n12134_o;
  assign n12136_o = {n11975_o, n12135_o};
  assign n12137_o = data_read[4:0];
  assign n12138_o = data_read[4:0];
  assign n12139_o = n12543_q[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n12140_o = n11922_o ? n12138_o : n12139_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n12141_o = n11925_o ? n12137_o : n12140_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1024:33  */
  assign n12142_o = n11956_o ? n12136_o : n12141_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1024:33  */
  assign n12143_o = n11956_o ? n11957_o : last_flags1;
  assign n12144_o = n12142_o[3:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1014:33  */
  assign n12145_o = z_error ? n11954_o : n12144_o;
  assign n12146_o = n12142_o[4];
  assign n12147_o = data_read[4];
  assign n12148_o = data_read[4];
  assign n12149_o = n12543_q[4];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n12150_o = n11922_o ? n12148_o : n12149_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n12151_o = n11925_o ? n12147_o : n12150_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1014:33  */
  assign n12152_o = z_error ? n12151_o : n12146_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1014:33  */
  assign n12153_o = z_error ? last_flags1 : n12143_o;
  assign n12154_o = {n12152_o, n12145_o};
  assign n12155_o = ccrin[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1012:33  */
  assign n12156_o = n11936_o ? n12155_o : n12154_o;
  assign n12157_o = ccrin[7:5];
  assign n12158_o = data_read[7:5];
  assign n12159_o = data_read[7:5];
  assign n12160_o = n12543_q[7:5];
  /* ../TG68K.C/TG68K_ALU.vhd:1000:33  */
  assign n12161_o = n11922_o ? n12159_o : n12160_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1003:33  */
  assign n12162_o = n11925_o ? n12158_o : n12161_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1012:33  */
  assign n12163_o = n11936_o ? n12157_o : n12162_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1012:33  */
  assign n12169_o = n11936_o ? last_flags1 : n12153_o;
  assign n12170_o = {n12163_o, n12156_o};
  /* ../TG68K.C/TG68K_ALU.vhd:999:25  */
  assign n12172_o = clkena_lw ? n12169_o : last_flags1;
  /* ../TG68K.C/TG68K_ALU.vhd:999:25  */
  assign n12173_o = clkena_lw ? n11935_o : asl_vflag;
  /* ../TG68K.C/TG68K_ALU.vhd:997:25  */
  assign n12176_o = reset ? last_flags1 : n12172_o;
  /* ../TG68K.C/TG68K_ALU.vhd:997:25  */
  assign n12177_o = reset ? asl_vflag : n12173_o;
  assign n12179_o = n12174_o[4:0];
  assign n12180_o = n12170_o[4:0];
  assign n12181_o = n12543_q[4:0];
  /* ../TG68K.C/TG68K_ALU.vhd:999:25  */
  assign n12182_o = clkena_lw ? n12180_o : n12181_o;
  /* ../TG68K.C/TG68K_ALU.vhd:997:25  */
  assign n12183_o = reset ? n12179_o : n12182_o;
  assign n12184_o = {3'b000, n12183_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1128:38  */
  assign n12191_o = exe_opcode[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1129:59  */
  assign n12192_o = reg_qa[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1129:49  */
  assign n12193_o = signedop & n12192_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1129:33  */
  assign n12196_o = n12193_o ? 32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:1134:59  */
  assign n12197_o = op2out[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1134:49  */
  assign n12198_o = signedop & n12197_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1134:33  */
  assign n12201_o = n12198_o ? 32'b11111111111111111111111111111111 : 32'b00000000000000000000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:1140:63  */
  assign n12202_o = reg_qa[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1141:63  */
  assign n12203_o = op2out[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1142:59  */
  assign n12204_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1142:49  */
  assign n12205_o = signedop & n12204_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1142:33  */
  assign n12208_o = n12205_o ? 16'b1111111111111111 : 16'b0000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:1147:59  */
  assign n12209_o = op2out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1147:49  */
  assign n12210_o = signedop & n12209_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1147:33  */
  assign n12213_o = n12210_o ? 16'b1111111111111111 : 16'b0000000000000000;
  assign n12214_o = {n12208_o, n12202_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1128:25  */
  assign n12215_o = n12191_o ? n12196_o : n12214_o;
  assign n12216_o = {n12213_o, n12203_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1128:25  */
  assign n12217_o = n12191_o ? n12201_o : n12216_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1153:62  */
  assign n12218_o = faktora[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1153:77  */
  assign n12219_o = {n12218_o, faktora};
  /* ../TG68K.C/TG68K_ALU.vhd:1153:108  */
  assign n12220_o = reg_qa[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1153:100  */
  assign n12221_o = {n12219_o, n12220_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1153:133  */
  assign n12222_o = faktorb[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1153:148  */
  assign n12223_o = {n12222_o, faktorb};
  /* ../TG68K.C/TG68K_ALU.vhd:1153:179  */
  assign n12224_o = op2out[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1153:171  */
  assign n12225_o = {n12223_o, n12224_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1153:123  */
  assign n12226_o = {64'b0, n12221_o};  //  uext
  /* ../TG68K.C/TG68K_ALU.vhd:1153:123  */
  assign n12227_o = {64'b0, n12225_o};  //  uext
  /* ../TG68K.C/TG68K_ALU.vhd:1153:123  */
  assign n12228_o = n12226_o * n12227_o; // umul
  /* ../TG68K.C/TG68K_ALU.vhd:1201:32  */
  assign n12229_o = result_mulu[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:1201:46  */
  assign n12231_o = n12229_o == 32'b00000000000000000000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:1201:72  */
  assign n12232_o = ~signedop;
  /* ../TG68K.C/TG68K_ALU.vhd:1201:91  */
  assign n12233_o = result_mulu[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1201:95  */
  assign n12234_o = ~n12233_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1201:77  */
  assign n12235_o = n12232_o | n12234_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1201:59  */
  assign n12236_o = n12231_o & n12235_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1202:37  */
  assign n12237_o = result_mulu[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:1202:51  */
  assign n12239_o = n12237_o == 32'b11111111111111111111111111111111;
  /* ../TG68K.C/TG68K_ALU.vhd:1202:64  */
  assign n12240_o = n12239_o & signedop;
  /* ../TG68K.C/TG68K_ALU.vhd:1202:96  */
  assign n12241_o = result_mulu[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1202:81  */
  assign n12242_o = n12240_o & n12241_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1201:102  */
  assign n12243_o = n12236_o | n12242_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1201:17  */
  assign n12246_o = n12243_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:1227:77  */
  assign n12251_o = result_mulu[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:1240:32  */
  assign n12259_o = opcode[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1240:47  */
  assign n12260_o = opcode[8];
  /* ../TG68K.C/TG68K_ALU.vhd:1240:37  */
  assign n12261_o = n12259_o & n12260_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1240:66  */
  assign n12262_o = opcode[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1240:56  */
  assign n12263_o = ~n12262_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1240:81  */
  assign n12264_o = sndopc[11];
  /* ../TG68K.C/TG68K_ALU.vhd:1240:71  */
  assign n12265_o = n12263_o & n12264_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1240:52  */
  assign n12266_o = n12261_o | n12265_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12268_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12269_o = divs & n12268_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12270_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12271_o = divs & n12270_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12272_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12273_o = divs & n12272_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12274_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12275_o = divs & n12274_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12276_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12277_o = divs & n12276_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12278_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12279_o = divs & n12278_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12280_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12281_o = divs & n12280_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12282_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12283_o = divs & n12282_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12284_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12285_o = divs & n12284_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12286_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12287_o = divs & n12286_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12288_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12289_o = divs & n12288_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12290_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12291_o = divs & n12290_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12292_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12293_o = divs & n12292_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12294_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12295_o = divs & n12294_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12296_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12297_o = divs & n12296_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12298_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12299_o = divs & n12298_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12300_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12301_o = divs & n12300_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12302_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12303_o = divs & n12302_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12304_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12305_o = divs & n12304_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12306_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12307_o = divs & n12306_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12308_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12309_o = divs & n12308_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12310_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12311_o = divs & n12310_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12312_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12313_o = divs & n12312_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12314_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12315_o = divs & n12314_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12316_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12317_o = divs & n12316_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12318_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12319_o = divs & n12318_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12320_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12321_o = divs & n12320_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12322_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12323_o = divs & n12322_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12324_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12325_o = divs & n12324_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12326_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12327_o = divs & n12326_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12328_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12329_o = divs & n12328_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1242:68  */
  assign n12330_o = reg_qa[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1242:58  */
  assign n12331_o = divs & n12330_o;
  assign n12332_o = {n12269_o, n12271_o, n12273_o, n12275_o};
  assign n12333_o = {n12277_o, n12279_o, n12281_o, n12283_o};
  assign n12334_o = {n12285_o, n12287_o, n12289_o, n12291_o};
  assign n12335_o = {n12293_o, n12295_o, n12297_o, n12299_o};
  assign n12336_o = {n12301_o, n12303_o, n12305_o, n12307_o};
  assign n12337_o = {n12309_o, n12311_o, n12313_o, n12315_o};
  assign n12338_o = {n12317_o, n12319_o, n12321_o, n12323_o};
  assign n12339_o = {n12325_o, n12327_o, n12329_o, n12331_o};
  assign n12340_o = {n12332_o, n12333_o, n12334_o, n12335_o};
  assign n12341_o = {n12336_o, n12337_o, n12338_o, n12339_o};
  assign n12342_o = {n12340_o, n12341_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1243:30  */
  assign n12343_o = exe_opcode[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1243:39  */
  assign n12345_o = n12343_o | 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:1245:52  */
  assign n12346_o = result_div_pre[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1248:38  */
  assign n12347_o = exe_opcode[14];
  /* ../TG68K.C/TG68K_ALU.vhd:1248:57  */
  assign n12348_o = sndopc[10];
  /* ../TG68K.C/TG68K_ALU.vhd:1248:47  */
  assign n12349_o = n12347_o & n12348_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1248:25  */
  assign n12350_o = n12349_o ? reg_qb : n12342_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1251:52  */
  assign n12351_o = result_div_pre[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1243:17  */
  assign n12352_o = n12345_o ? n12346_o : n12351_o;
  assign n12353_o = {n12350_o, reg_qa};
  assign n12354_o = n12353_o[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1243:17  */
  assign n12355_o = n12345_o ? 16'b0000000000000000 : n12354_o;
  assign n12356_o = n12353_o[47:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1243:17  */
  assign n12357_o = n12345_o ? reg_qa : n12356_o;
  assign n12358_o = n12353_o[63:48];
  assign n12359_o = n12342_o[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1243:17  */
  assign n12360_o = n12345_o ? n12359_o : n12358_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1253:42  */
  assign n12362_o = opcode[15];
  /* ../TG68K.C/TG68K_ALU.vhd:1253:46  */
  assign n12363_o = ~n12362_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1253:33  */
  assign n12364_o = signedop | n12363_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1254:44  */
  assign n12365_o = op2out[31:16];
  /* ../TG68K.C/TG68K_ALU.vhd:1253:17  */
  assign n12367_o = n12364_o ? n12365_o : 16'b0000000000000000;
  /* ../TG68K.C/TG68K_ALU.vhd:1258:43  */
  assign n12368_o = op2out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1258:33  */
  assign n12369_o = signedop & n12368_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1259:44  */
  assign n12370_o = div_reg[63:31];
  /* ../TG68K.C/TG68K_ALU.vhd:1259:64  */
  assign n12372_o = {1'b1, op2out};
  /* ../TG68K.C/TG68K_ALU.vhd:1259:59  */
  assign n12373_o = n12370_o + n12372_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1261:44  */
  assign n12374_o = div_reg[63:31];
  /* ../TG68K.C/TG68K_ALU.vhd:1261:64  */
  assign n12376_o = {1'b0, op2outext};
  /* ../TG68K.C/TG68K_ALU.vhd:1261:94  */
  assign n12377_o = op2out[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1261:87  */
  assign n12378_o = {n12376_o, n12377_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1261:59  */
  assign n12379_o = n12374_o - n12378_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1258:17  */
  assign n12380_o = n12369_o ? n12373_o : n12379_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1266:43  */
  assign n12381_o = div_sub[32];
  /* ../TG68K.C/TG68K_ALU.vhd:1269:58  */
  assign n12382_o = div_reg[62:31];
  /* ../TG68K.C/TG68K_ALU.vhd:1271:58  */
  assign n12383_o = div_sub[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1268:17  */
  assign n12384_o = div_bit ? n12382_o : n12383_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1273:49  */
  assign n12385_o = div_reg[30:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1273:63  */
  assign n12386_o = ~div_bit;
  /* ../TG68K.C/TG68K_ALU.vhd:1273:62  */
  assign n12387_o = {n12385_o, n12386_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1276:66  */
  assign n12388_o = div_quot[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1276:57  */
  assign n12390_o = 32'b00000000000000000000000000000000 - n12388_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1279:64  */
  assign n12391_o = div_quot[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1275:17  */
  assign n12392_o = div_neg ? n12390_o : n12391_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1282:44  */
  assign n12393_o = ~div_bit;
  /* ../TG68K.C/TG68K_ALU.vhd:1282:34  */
  assign n12394_o = nozero | n12393_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1282:50  */
  assign n12395_o = n12394_o & signedop;
  /* ../TG68K.C/TG68K_ALU.vhd:1282:78  */
  assign n12396_o = op2out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1282:83  */
  assign n12397_o = n12396_o ^ op1_sign;
  /* ../TG68K.C/TG68K_ALU.vhd:1282:96  */
  assign n12398_o = n12397_o ^ div_qsign;
  /* ../TG68K.C/TG68K_ALU.vhd:1282:67  */
  assign n12399_o = n12395_o & n12398_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1283:37  */
  assign n12400_o = ~signedop;
  /* ../TG68K.C/TG68K_ALU.vhd:1283:54  */
  assign n12401_o = div_over[32];
  /* ../TG68K.C/TG68K_ALU.vhd:1283:58  */
  assign n12402_o = ~n12401_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1283:42  */
  assign n12403_o = n12400_o & n12402_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1283:25  */
  assign n12404_o = n12399_o | n12403_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1283:65  */
  assign n12406_o = n12404_o & 1'b1;
  /* ../TG68K.C/TG68K_ALU.vhd:1282:17  */
  assign n12409_o = n12406_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:1294:47  */
  assign n12415_o = micro_state != 7'b1011010;
  /* ../TG68K.C/TG68K_ALU.vhd:1298:47  */
  assign n12418_o = micro_state == 7'b1010101;
  /* ../TG68K.C/TG68K_ALU.vhd:1300:65  */
  assign n12419_o = dividend[63];
  /* ../TG68K.C/TG68K_ALU.vhd:1300:53  */
  assign n12420_o = divs & n12419_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1302:61  */
  assign n12422_o = 64'b0000000000000000000000000000000000000000000000000000000000000000 - dividend;
  /* ../TG68K.C/TG68K_ALU.vhd:1300:41  */
  assign n12423_o = n12420_o ? n12422_o : dividend;
  /* ../TG68K.C/TG68K_ALU.vhd:1300:41  */
  assign n12426_o = n12420_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68K_ALU.vhd:1309:51  */
  assign n12427_o = ~div_bit;
  /* ../TG68K.C/TG68K_ALU.vhd:1309:63  */
  assign n12428_o = n12427_o | nozero;
  /* ../TG68K.C/TG68K_ALU.vhd:1298:33  */
  assign n12429_o = n12418_o ? n12423_o : div_quot;
  /* ../TG68K.C/TG68K_ALU.vhd:1298:33  */
  assign n12431_o = n12418_o ? 1'b0 : n12428_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1311:47  */
  assign n12434_o = micro_state == 7'b1010110;
  /* ../TG68K.C/TG68K_ALU.vhd:1312:72  */
  assign n12435_o = op2out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:1312:77  */
  assign n12436_o = n12435_o ^ op1_sign;
  /* ../TG68K.C/TG68K_ALU.vhd:1312:61  */
  assign n12437_o = signedop & n12436_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1316:73  */
  assign n12438_o = div_reg[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:1316:65  */
  assign n12440_o = {1'b0, n12438_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1316:93  */
  assign n12442_o = {1'b0, op2outext};
  /* ../TG68K.C/TG68K_ALU.vhd:1316:123  */
  assign n12443_o = op2out[15:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1316:116  */
  assign n12444_o = {n12442_o, n12443_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1316:88  */
  assign n12445_o = n12440_o - n12444_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1319:40  */
  assign n12448_o = exec[68];
  /* ../TG68K.C/TG68K_ALU.vhd:1319:56  */
  assign n12449_o = ~n12448_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1322:87  */
  assign n12450_o = div_quot[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:1322:78  */
  assign n12452_o = 32'b00000000000000000000000000000000 - n12450_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1324:85  */
  assign n12453_o = div_quot[63:32];
  /* ../TG68K.C/TG68K_ALU.vhd:1321:41  */
  assign n12454_o = op1_sign ? n12452_o : n12453_o;
  assign n12455_o = {n12454_o, result_div_pre};
  /* ../TG68K.C/TG68K_ALU.vhd:1293:25  */
  assign n12457_o = clkena_lw & n12449_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1293:25  */
  assign n12458_o = clkena_lw & n12415_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1293:25  */
  assign n12460_o = clkena_lw & n12434_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1293:25  */
  assign n12461_o = clkena_lw & n12434_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1293:25  */
  assign n12464_o = clkena_lw & n12418_o;
  assign n12474_o = {n9634_o, n9631_o};
  assign n12475_o = {n9785_o, n9778_o, n9771_o};
  assign n12476_o = {n9763_o, n9762_o, n9757_o, n9715_o};
  /* ../TG68K.C/TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12477_q <= n12176_o;
  /* ../TG68K.C/TG68K_ALU.vhd:996:17  */
  assign n12478_o = {n9807_o, n9845_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12479_o = n12457_o ? n12455_o : result_div;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12480_q <= n12479_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12481_o = n12458_o ? n12409_o : v_flag;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12482_q <= n12481_o;
  /* ../TG68K.C/TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12483_q <= n12177_o;
  /* ../TG68K.C/TG68K_ALU.vhd:405:17  */
  assign n12485_o = clkena_lw ? n9866_o : bchg;
  /* ../TG68K.C/TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n12486_q <= n12485_o;
  /* ../TG68K.C/TG68K_ALU.vhd:405:17  */
  assign n12487_o = clkena_lw ? n9870_o : bset;
  /* ../TG68K.C/TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n12488_q <= n12487_o;
  assign n12492_o = mulu_reg[31:0];
  /* ../TG68K.C/TG68K_ALU.vhd:1211:17  */
  assign n12493_o = clkena_lw ? n12251_o : n12492_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1211:17  */
  always @(posedge clk)
    n12494_q <= n12493_o;
  assign n12496_o = {32'bZ, n12494_q};
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12498_o = clkena_lw ? n12429_o : div_reg;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12499_q <= n12498_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12500_o = {n12384_o, n12387_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12502_o = n12460_o ? n12437_o : div_neg;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12503_q <= n12502_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12504_o = n12461_o ? n12445_o : div_over;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12505_q <= n12504_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12506_o = clkena_lw ? n12431_o : nozero;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12507_q <= n12506_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12508_o = {n12360_o, n12357_o, n12355_o};
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12509_o = clkena_lw ? divs : signedop;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12510_q <= n12509_o;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12511_o = n12464_o ? n12426_o : op1_sign;
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12512_q <= n12511_o;
  assign n12515_o = {n10445_o, n10433_o, n10418_o, n10403_o, n10388_o, n10373_o, n10358_o, n10343_o, n10328_o, n10313_o, n10298_o, n10283_o, n10268_o, n10253_o, n10238_o, n10223_o, n10208_o, n10193_o, n10178_o, n10163_o, n10148_o, n10133_o, n10118_o, n10103_o, n10088_o, n10073_o, n10058_o, n10043_o, n10028_o, n10013_o, n9998_o, n9982_o};
  assign n12517_o = {n11208_o, n11198_o, n11181_o, n11164_o, n11147_o, n11130_o, n11113_o, n11096_o, n11079_o, n11062_o, n11045_o, n11028_o, n11011_o, n10994_o, n10977_o, n10960_o, n10943_o, n10926_o, n10909_o, n10892_o, n10875_o, n10858_o, n10841_o, n10824_o, n10807_o, n10790_o, n10773_o, n10756_o, n10739_o, n10722_o, n10705_o, n10688_o, n10671_o, n10654_o, n10637_o, n10620_o, n10603_o, n10586_o, n10569_o, n10552_o};
  assign n12518_o = {n10446_o, n10438_o, n10423_o, n10408_o, n10393_o, n10378_o, n10363_o, n10348_o, n10333_o, n10318_o, n10303_o, n10288_o, n10273_o, n10258_o, n10243_o, n10228_o, n10213_o, n10198_o, n10183_o, n10168_o, n10153_o, n10138_o, n10123_o, n10108_o, n10093_o, n10078_o, n10063_o, n10048_o, n10033_o, n10018_o, n10003_o, n9987_o};
  assign n12520_o = {n10502_o, n10503_o};
  assign n12521_o = {n11292_o, n11321_o, n11318_o};
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12522_o = clkena_lw ? n9929_o : bf_bset;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12523_q <= n12522_o;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12524_o = clkena_lw ? n9933_o : bf_bchg;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12525_q <= n12524_o;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12526_o = clkena_lw ? n9937_o : bf_ins;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12527_q <= n12526_o;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12528_o = clkena_lw ? n9941_o : bf_exts;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12529_q <= n12528_o;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12530_o = clkena_lw ? n9945_o : bf_fffo;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12531_q <= n12530_o;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12532_o = clkena_lw ? n9954_o : bf_d32;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12533_q <= n12532_o;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12534_o = clkena_lw ? n9948_o : bf_s32;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12535_q <= n12534_o;
  assign n12537_o = {n11812_o, n11810_o, n11807_o, n11804_o, n11801_o, n11814_o};
  assign n12538_o = {n11493_o, n11490_o, n11494_o, n11488_o, n11492_o};
  assign n12539_o = {n11747_o, n11749_o};
  assign n12540_o = {n11828_o, n11823_o, n11834_o};
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12541_o = clkena_lw ? n9956_o : n12542_q;
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12542_q <= n12541_o;
  /* ../TG68K.C/TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12543_q <= n12184_o;
  /* ../TG68K.C/TG68K_ALU.vhd:76:17  */
  assign n12544_o = op1out[0];
  /* ../TG68K.C/TG68K_ALU.vhd:75:17  */
  assign n12545_o = op1out[1];
  /* ../TG68K.C/TG68K_ALU.vhd:74:17  */
  assign n12546_o = op1out[2];
  /* ../TG68K.C/TG68K_ALU.vhd:73:17  */
  assign n12547_o = op1out[3];
  /* ../TG68K.C/TG68K_ALU.vhd:72:17  */
  assign n12548_o = op1out[4];
  /* ../TG68K.C/TG68K_ALU.vhd:66:17  */
  assign n12549_o = op1out[5];
  /* ../TG68K.C/TG68K_ALU.vhd:446:17  */
  assign n12550_o = op1out[6];
  assign n12551_o = op1out[7];
  assign n12552_o = op1out[8];
  assign n12553_o = op1out[9];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12554_o = op1out[10];
  assign n12555_o = op1out[11];
  assign n12556_o = op1out[12];
  assign n12557_o = op1out[13];
  assign n12558_o = op1out[14];
  /* ../TG68K.C/TG68K_ALU.vhd:405:17  */
  assign n12559_o = op1out[15];
  /* ../TG68K.C/TG68K_ALU.vhd:996:17  */
  assign n12560_o = op1out[16];
  assign n12561_o = op1out[17];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12562_o = op1out[18];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12563_o = op1out[19];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12564_o = op1out[20];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12565_o = op1out[21];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12566_o = op1out[22];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12567_o = op1out[23];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12568_o = op1out[24];
  /* ../TG68K.C/TG68K_ALU.vhd:1292:17  */
  assign n12569_o = op1out[25];
  /* ../TG68K.C/TG68K_ALU.vhd:1290:1  */
  assign n12570_o = op1out[26];
  assign n12571_o = op1out[27];
  assign n12572_o = op1out[28];
  /* ../TG68K.C/TG68K_ALU.vhd:1237:1  */
  assign n12573_o = op1out[29];
  assign n12574_o = op1out[30];
  /* ../TG68K.C/TG68K_ALU.vhd:1211:17  */
  assign n12575_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12576_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12576_o)
      2'b00: n12577_o = n12544_o;
      2'b01: n12577_o = n12545_o;
      2'b10: n12577_o = n12546_o;
      2'b11: n12577_o = n12547_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12578_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12578_o)
      2'b00: n12579_o = n12548_o;
      2'b01: n12579_o = n12549_o;
      2'b10: n12579_o = n12550_o;
      2'b11: n12579_o = n12551_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12580_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12580_o)
      2'b00: n12581_o = n12552_o;
      2'b01: n12581_o = n12553_o;
      2'b10: n12581_o = n12554_o;
      2'b11: n12581_o = n12555_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12582_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12582_o)
      2'b00: n12583_o = n12556_o;
      2'b01: n12583_o = n12557_o;
      2'b10: n12583_o = n12558_o;
      2'b11: n12583_o = n12559_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12584_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12584_o)
      2'b00: n12585_o = n12560_o;
      2'b01: n12585_o = n12561_o;
      2'b10: n12585_o = n12562_o;
      2'b11: n12585_o = n12563_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12586_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12586_o)
      2'b00: n12587_o = n12564_o;
      2'b01: n12587_o = n12565_o;
      2'b10: n12587_o = n12566_o;
      2'b11: n12587_o = n12567_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12588_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12588_o)
      2'b00: n12589_o = n12568_o;
      2'b01: n12589_o = n12569_o;
      2'b10: n12589_o = n12570_o;
      2'b11: n12589_o = n12571_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12590_o = bit_number[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12590_o)
      2'b00: n12591_o = n12572_o;
      2'b01: n12591_o = n12573_o;
      2'b10: n12591_o = n12574_o;
      2'b11: n12591_o = n12575_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12592_o = bit_number[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12592_o)
      2'b00: n12593_o = n12577_o;
      2'b01: n12593_o = n12579_o;
      2'b10: n12593_o = n12581_o;
      2'b11: n12593_o = n12583_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12594_o = bit_number[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  always @*
    case (n12594_o)
      2'b00: n12595_o = n12585_o;
      2'b01: n12595_o = n12587_o;
      2'b10: n12595_o = n12589_o;
      2'b11: n12595_o = n12591_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12596_o = bit_number[4];
  /* ../TG68K.C/TG68K_ALU.vhd:433:37  */
  assign n12597_o = n12596_o ? n12595_o : n12593_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12598_o = bit_number[4];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12599_o = ~n12598_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12600_o = bit_number[3];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12601_o = ~n12600_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12602_o = n12599_o & n12601_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12603_o = n12599_o & n12600_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12604_o = n12598_o & n12601_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12605_o = n12598_o & n12600_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12606_o = bit_number[2];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12607_o = ~n12606_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12608_o = n12602_o & n12607_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12609_o = n12602_o & n12606_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12610_o = n12603_o & n12607_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12611_o = n12603_o & n12606_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12612_o = n12604_o & n12607_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12613_o = n12604_o & n12606_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12614_o = n12605_o & n12607_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12615_o = n12605_o & n12606_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12616_o = bit_number[1];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12617_o = ~n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12618_o = n12608_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12619_o = n12608_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12620_o = n12609_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12621_o = n12609_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12622_o = n12610_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12623_o = n12610_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12624_o = n12611_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12625_o = n12611_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12626_o = n12612_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12627_o = n12612_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12628_o = n12613_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12629_o = n12613_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12630_o = n12614_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12631_o = n12614_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12632_o = n12615_o & n12617_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12633_o = n12615_o & n12616_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12634_o = bit_number[0];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12635_o = ~n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12636_o = n12618_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12637_o = n12618_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12638_o = n12619_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12639_o = n12619_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12640_o = n12620_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12641_o = n12620_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12642_o = n12621_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12643_o = n12621_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12644_o = n12622_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12645_o = n12622_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12646_o = n12623_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12647_o = n12623_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12648_o = n12624_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12649_o = n12624_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12650_o = n12625_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12651_o = n12625_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12652_o = n12626_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12653_o = n12626_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12654_o = n12627_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12655_o = n12627_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12656_o = n12628_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12657_o = n12628_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12658_o = n12629_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12659_o = n12629_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12660_o = n12630_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12661_o = n12630_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12662_o = n12631_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12663_o = n12631_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12664_o = n12632_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12665_o = n12632_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12666_o = n12633_o & n12635_o;
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12667_o = n12633_o & n12634_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12668_o = op1out[0];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12669_o = n12636_o ? n9902_o : n12668_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12670_o = op1out[1];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12671_o = n12637_o ? n9902_o : n12670_o;
  assign n12672_o = op1out[2];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12673_o = n12638_o ? n9902_o : n12672_o;
  assign n12674_o = op1out[3];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12675_o = n12639_o ? n9902_o : n12674_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12676_o = op1out[4];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12677_o = n12640_o ? n9902_o : n12676_o;
  assign n12678_o = op1out[5];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12679_o = n12641_o ? n9902_o : n12678_o;
  assign n12680_o = op1out[6];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12681_o = n12642_o ? n9902_o : n12680_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12682_o = op1out[7];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12683_o = n12643_o ? n9902_o : n12682_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12684_o = op1out[8];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12685_o = n12644_o ? n9902_o : n12684_o;
  assign n12686_o = op1out[9];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12687_o = n12645_o ? n9902_o : n12686_o;
  assign n12688_o = op1out[10];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12689_o = n12646_o ? n9902_o : n12688_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12690_o = op1out[11];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12691_o = n12647_o ? n9902_o : n12690_o;
  assign n12692_o = op1out[12];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12693_o = n12648_o ? n9902_o : n12692_o;
  assign n12694_o = op1out[13];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12695_o = n12649_o ? n9902_o : n12694_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12696_o = op1out[14];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12697_o = n12650_o ? n9902_o : n12696_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12698_o = op1out[15];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12699_o = n12651_o ? n9902_o : n12698_o;
  assign n12700_o = op1out[16];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12701_o = n12652_o ? n9902_o : n12700_o;
  assign n12702_o = op1out[17];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12703_o = n12653_o ? n9902_o : n12702_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12704_o = op1out[18];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12705_o = n12654_o ? n9902_o : n12704_o;
  assign n12706_o = op1out[19];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12707_o = n12655_o ? n9902_o : n12706_o;
  assign n12708_o = op1out[20];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12709_o = n12656_o ? n9902_o : n12708_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12710_o = op1out[21];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12711_o = n12657_o ? n9902_o : n12710_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12712_o = op1out[22];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12713_o = n12658_o ? n9902_o : n12712_o;
  assign n12714_o = op1out[23];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12715_o = n12659_o ? n9902_o : n12714_o;
  assign n12716_o = op1out[24];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12717_o = n12660_o ? n9902_o : n12716_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12718_o = op1out[25];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12719_o = n12661_o ? n9902_o : n12718_o;
  assign n12720_o = op1out[26];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12721_o = n12662_o ? n9902_o : n12720_o;
  assign n12722_o = op1out[27];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12723_o = n12663_o ? n9902_o : n12722_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12724_o = op1out[28];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12725_o = n12664_o ? n9902_o : n12724_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12726_o = op1out[29];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12727_o = n12665_o ? n9902_o : n12726_o;
  assign n12728_o = op1out[30];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12729_o = n12666_o ? n9902_o : n12728_o;
  assign n12730_o = op1out[31];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12731_o = n12667_o ? n9902_o : n12730_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12732_o = {n12731_o, n12729_o, n12727_o, n12725_o, n12723_o, n12721_o, n12719_o, n12717_o, n12715_o, n12713_o, n12711_o, n12709_o, n12707_o, n12705_o, n12703_o, n12701_o, n12699_o, n12697_o, n12695_o, n12693_o, n12691_o, n12689_o, n12687_o, n12685_o, n12683_o, n12681_o, n12679_o, n12677_o, n12675_o, n12673_o, n12671_o, n12669_o};
  /* ../TG68K.C/TG68K_ALU.vhd:435:26  */
  assign n12733_o = datareg[0];
  /* ../TG68K.C/TG68K_ALU.vhd:435:17  */
  assign n12734_o = datareg[1];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12735_o = datareg[2];
  assign n12736_o = datareg[3];
  assign n12737_o = datareg[4];
  assign n12738_o = datareg[5];
  assign n12739_o = datareg[6];
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12740_o = datareg[7];
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12741_o = datareg[8];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12742_o = datareg[9];
  assign n12743_o = datareg[10];
  assign n12744_o = datareg[11];
  assign n12745_o = datareg[12];
  assign n12746_o = datareg[13];
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12747_o = datareg[14];
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12748_o = datareg[15];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12749_o = datareg[16];
  assign n12750_o = datareg[17];
  assign n12751_o = datareg[18];
  assign n12752_o = datareg[19];
  assign n12753_o = datareg[20];
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12754_o = datareg[21];
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12755_o = datareg[22];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12756_o = datareg[23];
  assign n12757_o = datareg[24];
  assign n12758_o = datareg[25];
  assign n12759_o = datareg[26];
  assign n12760_o = datareg[27];
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12761_o = datareg[28];
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12762_o = datareg[29];
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12763_o = datareg[30];
  assign n12764_o = datareg[31];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12765_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12765_o)
      2'b00: n12766_o = n12733_o;
      2'b01: n12766_o = n12734_o;
      2'b10: n12766_o = n12735_o;
      2'b11: n12766_o = n12736_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12767_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12767_o)
      2'b00: n12768_o = n12737_o;
      2'b01: n12768_o = n12738_o;
      2'b10: n12768_o = n12739_o;
      2'b11: n12768_o = n12740_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12769_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12769_o)
      2'b00: n12770_o = n12741_o;
      2'b01: n12770_o = n12742_o;
      2'b10: n12770_o = n12743_o;
      2'b11: n12770_o = n12744_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12771_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12771_o)
      2'b00: n12772_o = n12745_o;
      2'b01: n12772_o = n12746_o;
      2'b10: n12772_o = n12747_o;
      2'b11: n12772_o = n12748_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12773_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12773_o)
      2'b00: n12774_o = n12749_o;
      2'b01: n12774_o = n12750_o;
      2'b10: n12774_o = n12751_o;
      2'b11: n12774_o = n12752_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12775_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12775_o)
      2'b00: n12776_o = n12753_o;
      2'b01: n12776_o = n12754_o;
      2'b10: n12776_o = n12755_o;
      2'b11: n12776_o = n12756_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12777_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12777_o)
      2'b00: n12778_o = n12757_o;
      2'b01: n12778_o = n12758_o;
      2'b10: n12778_o = n12759_o;
      2'b11: n12778_o = n12760_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12779_o = n10448_o[1:0];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12779_o)
      2'b00: n12780_o = n12761_o;
      2'b01: n12780_o = n12762_o;
      2'b10: n12780_o = n12763_o;
      2'b11: n12780_o = n12764_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12781_o = n10448_o[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12781_o)
      2'b00: n12782_o = n12766_o;
      2'b01: n12782_o = n12768_o;
      2'b10: n12782_o = n12770_o;
      2'b11: n12782_o = n12772_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12783_o = n10448_o[3:2];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  always @*
    case (n12783_o)
      2'b00: n12784_o = n12774_o;
      2'b01: n12784_o = n12776_o;
      2'b10: n12784_o = n12778_o;
      2'b11: n12784_o = n12780_o;
    endcase
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12785_o = n10448_o[4];
  /* ../TG68K.C/TG68K_ALU.vhd:496:36  */
  assign n12786_o = n12785_o ? n12784_o : n12782_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12787_o = bit_msb[5];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12788_o = ~n12787_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12789_o = bit_msb[4];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12790_o = ~n12789_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12791_o = n12788_o & n12790_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12792_o = n12788_o & n12789_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12793_o = n12787_o & n12790_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12794_o = bit_msb[3];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12795_o = ~n12794_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12796_o = n12791_o & n12795_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12797_o = n12791_o & n12794_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12798_o = n12792_o & n12795_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12799_o = n12792_o & n12794_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12800_o = n12793_o & n12795_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12801_o = bit_msb[2];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12802_o = ~n12801_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12803_o = n12796_o & n12802_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12804_o = n12796_o & n12801_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12805_o = n12797_o & n12802_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12806_o = n12797_o & n12801_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12807_o = n12798_o & n12802_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12808_o = n12798_o & n12801_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12809_o = n12799_o & n12802_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12810_o = n12799_o & n12801_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12811_o = n12800_o & n12802_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12812_o = bit_msb[1];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12813_o = ~n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12814_o = n12803_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12815_o = n12803_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12816_o = n12804_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12817_o = n12804_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12818_o = n12805_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12819_o = n12805_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12820_o = n12806_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12821_o = n12806_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12822_o = n12807_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12823_o = n12807_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12824_o = n12808_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12825_o = n12808_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12826_o = n12809_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12827_o = n12809_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12828_o = n12810_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12829_o = n12810_o & n12812_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12830_o = n12811_o & n12813_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12831_o = bit_msb[0];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12832_o = ~n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12833_o = n12814_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12834_o = n12814_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12835_o = n12815_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12836_o = n12815_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12837_o = n12816_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12838_o = n12816_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12839_o = n12817_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12840_o = n12817_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12841_o = n12818_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12842_o = n12818_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12843_o = n12819_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12844_o = n12819_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12845_o = n12820_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12846_o = n12820_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12847_o = n12821_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12848_o = n12821_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12849_o = n12822_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12850_o = n12822_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12851_o = n12823_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12852_o = n12823_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12853_o = n12824_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12854_o = n12824_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12855_o = n12825_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12856_o = n12825_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12857_o = n12826_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12858_o = n12826_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12859_o = n12827_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12860_o = n12827_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12861_o = n12828_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12862_o = n12828_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12863_o = n12829_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12864_o = n12829_o & n12831_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12865_o = n12830_o & n12832_o;
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12866_o = n12830_o & n12831_o;
  assign n12867_o = n11459_o[0];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12868_o = n12833_o ? 1'b1 : n12867_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12869_o = n11459_o[1];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12870_o = n12834_o ? 1'b1 : n12869_o;
  assign n12871_o = n11459_o[2];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12872_o = n12835_o ? 1'b1 : n12871_o;
  assign n12873_o = n11459_o[3];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12874_o = n12836_o ? 1'b1 : n12873_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12875_o = n11459_o[4];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12876_o = n12837_o ? 1'b1 : n12875_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12877_o = n11459_o[5];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12878_o = n12838_o ? 1'b1 : n12877_o;
  assign n12879_o = n11459_o[6];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12880_o = n12839_o ? 1'b1 : n12879_o;
  assign n12881_o = n11459_o[7];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12882_o = n12840_o ? 1'b1 : n12881_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12883_o = n11459_o[8];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12884_o = n12841_o ? 1'b1 : n12883_o;
  assign n12885_o = n11459_o[9];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12886_o = n12842_o ? 1'b1 : n12885_o;
  assign n12887_o = n11459_o[10];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12888_o = n12843_o ? 1'b1 : n12887_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12889_o = n11459_o[11];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12890_o = n12844_o ? 1'b1 : n12889_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12891_o = n11459_o[12];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12892_o = n12845_o ? 1'b1 : n12891_o;
  assign n12893_o = n11459_o[13];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12894_o = n12846_o ? 1'b1 : n12893_o;
  assign n12895_o = n11459_o[14];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12896_o = n12847_o ? 1'b1 : n12895_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12897_o = n11459_o[15];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12898_o = n12848_o ? 1'b1 : n12897_o;
  assign n12899_o = n11459_o[16];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12900_o = n12849_o ? 1'b1 : n12899_o;
  assign n12901_o = n11459_o[17];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12902_o = n12850_o ? 1'b1 : n12901_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12903_o = n11459_o[18];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12904_o = n12851_o ? 1'b1 : n12903_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12905_o = n11459_o[19];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12906_o = n12852_o ? 1'b1 : n12905_o;
  assign n12907_o = n11459_o[20];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12908_o = n12853_o ? 1'b1 : n12907_o;
  assign n12909_o = n11459_o[21];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12910_o = n12854_o ? 1'b1 : n12909_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12911_o = n11459_o[22];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12912_o = n12855_o ? 1'b1 : n12911_o;
  assign n12913_o = n11459_o[23];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12914_o = n12856_o ? 1'b1 : n12913_o;
  assign n12915_o = n11459_o[24];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12916_o = n12857_o ? 1'b1 : n12915_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12917_o = n11459_o[25];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12918_o = n12858_o ? 1'b1 : n12917_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12919_o = n11459_o[26];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12920_o = n12859_o ? 1'b1 : n12919_o;
  assign n12921_o = n11459_o[27];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12922_o = n12860_o ? 1'b1 : n12921_o;
  assign n12923_o = n11459_o[28];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12924_o = n12861_o ? 1'b1 : n12923_o;
  /* ../TG68K.C/TG68K_ALU.vhd:572:17  */
  assign n12925_o = n11459_o[29];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12926_o = n12862_o ? 1'b1 : n12925_o;
  assign n12927_o = n11459_o[30];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12928_o = n12863_o ? 1'b1 : n12927_o;
  assign n12929_o = n11459_o[31];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12930_o = n12864_o ? 1'b1 : n12929_o;
  /* ../TG68K.C/TG68K_ALU.vhd:581:17  */
  assign n12931_o = n11459_o[32];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12932_o = n12865_o ? 1'b1 : n12931_o;
  /* ../TG68K.C/TG68K_ALU.vhd:575:17  */
  assign n12933_o = n11459_o[33];
  /* ../TG68K.C/TG68K_ALU.vhd:761:17  */
  assign n12934_o = n12866_o ? 1'b1 : n12933_o;
  assign n12935_o = {n12934_o, n12932_o, n12930_o, n12928_o, n12926_o, n12924_o, n12922_o, n12920_o, n12918_o, n12916_o, n12914_o, n12912_o, n12910_o, n12908_o, n12906_o, n12904_o, n12902_o, n12900_o, n12898_o, n12896_o, n12894_o, n12892_o, n12890_o, n12888_o, n12886_o, n12884_o, n12882_o, n12880_o, n12878_o, n12876_o, n12874_o, n12872_o, n12870_o, n12868_o};
endmodule

module TG68KdotC_Kernel
  (input  clk,
   input  nreset,
   input  clkena_in,
   input  [15:0] data_in,
   input  [2:0] ipl,
   input  ipl_autovector,
   input  berr,
   input  [1:0] cpu,
   output [31:0] addr_out,
   output [15:0] data_write,
   output nwr,
   output nuds,
   output nlds,
   output [1:0] busstate,
   output longword,
   output nresetout,
   output [2:0] fc,
   output clr_berr,
   output skipFetch,
   output [31:0] regin_out,
   output [3:0] cacr_out,
   output [31:0] vbr_out);
  wire use_vbr_stackframe;
  wire [3:0] syncreset;
  wire reset;
  wire clkena_lw;
  wire [31:0] tg68_pc;
  wire [31:0] tmp_tg68_pc;
  wire [31:0] tg68_pc_add;
  wire [31:0] pc_dataa;
  wire [31:0] pc_datab;
  wire [31:0] memaddr;
  wire [1:0] state;
  wire [1:0] datatype;
  wire [1:0] set_datatype;
  wire [1:0] exe_datatype;
  wire [1:0] setstate;
  wire setaddrvalue;
  wire addrvalue;
  wire [15:0] opcode;
  wire [15:0] exe_opcode;
  wire [15:0] sndopc;
  wire [31:0] exe_pc;
  wire [31:0] last_opc_pc;
  wire [15:0] last_opc_read;
  wire [31:0] reg_qa;
  wire [31:0] reg_qb;
  wire wwrena;
  wire lwrena;
  wire bwrena;
  wire regwrena_now;
  wire [3:0] rf_dest_addr;
  wire [3:0] rf_source_addr;
  wire [3:0] rf_source_addrd;
  wire [31:0] regin;
  wire [3:0] rdindex_a;
  wire [3:0] rdindex_b;
  wire wr_areg;
  wire [31:0] addr;
  wire [31:0] memaddr_reg;
  wire [31:0] memaddr_delta;
  wire [31:0] memaddr_delta_rega;
  wire [31:0] memaddr_delta_regb;
  wire use_base;
  wire [31:0] ea_data;
  wire [31:0] op1out;
  wire [31:0] op2out;
  wire [15:0] op1outbrief;
  wire [31:0] aluout;
  wire [31:0] data_write_tmp;
  wire [31:0] data_write_muxin;
  wire [47:0] data_write_mux;
  wire nextpass;
  wire setnextpass;
  wire setdispbyte;
  wire setdisp;
  wire regdirectsource;
  wire [31:0] addsub_q;
  wire [31:0] briefdata;
  wire [2:0] c_out;
  wire [31:0] memaddr_a;
  wire tg68_pc_brw;
  wire tg68_pc_word;
  wire getbrief;
  wire [15:0] brief;
  wire data_is_source;
  wire store_in_tmp;
  wire write_back;
  wire exec_write_back;
  wire setstackaddr;
  wire writepc;
  wire writepcbig;
  wire set_writepcbig;
  wire writepcnext;
  wire setopcode;
  wire decodeopc;
  wire execopc;
  wire execopc_alu;
  wire setexecopc;
  wire endopc;
  wire setendopc;
  wire [7:0] flags;
  wire [7:0] flagssr;
  wire [7:0] srin;
  wire exec_direct;
  wire exec_tas;
  wire set_exec_tas;
  wire exe_condition;
  wire ea_only;
  wire source_areg;
  wire source_lowbits;
  wire source_ldrlbits;
  wire source_ldrmbits;
  wire source_2ndhbits;
  wire source_2ndmbits;
  wire source_2ndlbits;
  wire dest_areg;
  wire dest_ldrareg;
  wire dest_ldrhbits;
  wire dest_ldrlbits;
  wire dest_2ndhbits;
  wire dest_2ndlbits;
  wire dest_hbits;
  wire [1:0] rot_bits;
  wire [1:0] set_rot_bits;
  wire [5:0] rot_cnt;
  wire [5:0] set_rot_cnt;
  wire movem_actiond;
  wire [3:0] movem_regaddr;
  wire [3:0] movem_mux;
  wire movem_presub;
  wire movem_run;
  wire set_direct_data;
  wire use_direct_data;
  wire direct_data;
  wire set_v_flag;
  wire set_vectoraddr;
  wire writesr;
  wire trap_berr;
  wire trap_illegal;
  wire trap_addr_error;
  wire trap_priv;
  wire trap_trace;
  wire trap_1010;
  wire trap_1111;
  wire trap_trap;
  wire trap_trapv;
  wire trap_interrupt;
  wire trapmake;
  wire trapd;
  wire [7:0] trap_sr;
  wire make_trace;
  wire make_berr;
  wire usestackframe2;
  wire set_stop;
  wire stop;
  wire [31:0] trap_vector;
  wire [31:0] trap_vector_vbr;
  wire [31:0] usp;
  wire [2:0] ipl_nr;
  wire [2:0] ripl_nr;
  wire [7:0] ipl_vec;
  wire interrupt;
  wire setinterrupt;
  wire svmode;
  wire presvmode;
  wire suppress_base;
  wire set_suppress_base;
  wire set_z_error;
  wire z_error;
  wire ea_build_now;
  wire build_logical;
  wire build_bcd;
  wire [31:0] data_read;
  wire [7:0] bf_ext_in;
  wire [7:0] bf_ext_out;
  wire long_start;
  wire long_start_alu;
  wire non_aligned;
  wire check_aligned;
  wire long_done;
  wire [5:0] memmask;
  wire [5:0] set_memmask;
  wire [3:0] memread;
  wire [5:0] wbmemmask;
  wire [5:0] memmaskmux;
  wire oddout;
  wire set_oddout;
  wire pcbase;
  wire set_pcbase;
  wire [31:0] last_data_read;
  wire [31:0] last_data_in;
  wire [5:0] bf_offset;
  wire [5:0] bf_width;
  wire [5:0] bf_bhits;
  wire [5:0] bf_shift;
  wire [5:0] alu_width;
  wire [5:0] alu_bf_shift;
  wire [5:0] bf_loffset;
  wire [31:0] bf_full_offset;
  wire [31:0] alu_bf_ffo_offset;
  wire [5:0] alu_bf_loffset;
  wire [31:0] movec_data;
  wire [31:0] vbr;
  wire [3:0] cacr;
  wire [2:0] dfc;
  wire [2:0] sfc;
  wire [88:0] set;
  wire [88:0] set_exec;
  wire [88:0] exec;
  wire [6:0] micro_state;
  wire [6:0] next_micro_state;
  wire [15:0] n15_o;
  wire [15:0] n16_o;
  wire [7:0] alu_n17;
  wire [4:0] n18_o;
  wire alu_n19;
  wire [7:0] alu_n20;
  wire [2:0] alu_n21;
  wire [31:0] alu_n22;
  wire [31:0] alu_n23;
  wire [7:0] alu_bf_ext_out;
  wire alu_set_v_flag;
  wire [7:0] alu_flags;
  wire [2:0] alu_c_out;
  wire [31:0] alu_addsub_q;
  wire [31:0] alu_aluout;
  wire n36_o;
  wire n37_o;
  wire n38_o;
  wire n39_o;
  wire n40_o;
  wire n41_o;
  wire [1:0] n44_o;
  wire n46_o;
  wire [1:0] n47_o;
  wire n49_o;
  wire n50_o;
  wire n53_o;
  wire n58_o;
  wire n59_o;
  wire n62_o;
  wire n63_o;
  wire n65_o;
  wire [5:0] n66_o;
  wire [4:0] n67_o;
  wire [5:0] n69_o;
  wire n70_o;
  wire n71_o;
  wire n73_o;
  wire n74_o;
  wire n75_o;
  wire n78_o;
  wire n79_o;
  wire n83_o;
  wire [2:0] n85_o;
  wire [3:0] n87_o;
  wire n88_o;
  wire n89_o;
  wire n99_o;
  wire n101_o;
  wire n103_o;
  wire n106_o;
  wire n111_o;
  wire n112_o;
  wire [15:0] n113_o;
  wire [31:0] n114_o;
  wire [23:0] n115_o;
  wire [7:0] n116_o;
  wire [31:0] n117_o;
  wire n119_o;
  wire [1:0] n120_o;
  wire n122_o;
  wire n123_o;
  wire n124_o;
  wire n125_o;
  wire n126_o;
  wire n127_o;
  wire n128_o;
  wire n129_o;
  wire n130_o;
  wire n131_o;
  wire n132_o;
  wire n133_o;
  wire n134_o;
  wire n135_o;
  wire n136_o;
  wire n137_o;
  wire n138_o;
  wire n139_o;
  wire n140_o;
  wire n141_o;
  wire [3:0] n142_o;
  wire [3:0] n143_o;
  wire [3:0] n144_o;
  wire [3:0] n145_o;
  wire [15:0] n146_o;
  wire [15:0] n147_o;
  wire [15:0] n148_o;
  wire [15:0] n149_o;
  wire [15:0] n150_o;
  wire [15:0] n151_o;
  wire [15:0] n152_o;
  wire [15:0] n153_o;
  wire n156_o;
  wire n157_o;
  wire n158_o;
  wire n159_o;
  wire [7:0] n160_o;
  wire [7:0] n161_o;
  wire [7:0] n162_o;
  wire n165_o;
  wire n166_o;
  wire n167_o;
  wire n168_o;
  wire n169_o;
  wire n170_o;
  wire n171_o;
  wire n172_o;
  wire n173_o;
  wire n174_o;
  wire n175_o;
  wire n176_o;
  wire n177_o;
  wire n178_o;
  wire n179_o;
  wire n180_o;
  wire n181_o;
  wire n182_o;
  wire n183_o;
  wire n184_o;
  wire n185_o;
  wire n186_o;
  wire n187_o;
  wire n188_o;
  wire n189_o;
  wire n190_o;
  wire n191_o;
  wire n192_o;
  wire [3:0] n193_o;
  wire [3:0] n194_o;
  wire [3:0] n195_o;
  wire [3:0] n196_o;
  wire [15:0] n197_o;
  wire [15:0] n198_o;
  wire [15:0] n199_o;
  wire [15:0] n200_o;
  wire [15:0] n201_o;
  wire [31:0] n202_o;
  wire [31:0] n203_o;
  wire [15:0] n204_o;
  wire [31:0] n205_o;
  wire n206_o;
  wire [31:0] n207_o;
  wire [31:0] n209_o;
  wire [31:0] n210_o;
  wire n214_o;
  wire n215_o;
  wire n216_o;
  wire n217_o;
  wire n221_o;
  wire [31:0] n222_o;
  wire n223_o;
  wire n224_o;
  wire [15:0] n226_o;
  wire [47:0] n227_o;
  wire [39:0] n228_o;
  wire [47:0] n230_o;
  wire [47:0] n231_o;
  wire n232_o;
  wire n233_o;
  wire [15:0] n234_o;
  wire n235_o;
  wire n236_o;
  wire [15:0] n237_o;
  wire [1:0] n238_o;
  wire n240_o;
  wire [7:0] n241_o;
  wire [7:0] n242_o;
  wire [15:0] n243_o;
  wire [1:0] n244_o;
  wire n246_o;
  wire [7:0] n247_o;
  wire [7:0] n248_o;
  wire [15:0] n249_o;
  wire [15:0] n250_o;
  wire [15:0] n251_o;
  wire [15:0] n252_o;
  wire [15:0] n253_o;
  wire [15:0] n254_o;
  wire n255_o;
  wire [7:0] n256_o;
  wire [7:0] n257_o;
  wire [15:0] n258_o;
  wire [15:0] n259_o;
  wire n272_o;
  wire n280_o;
  wire n283_o;
  wire n287_o;
  wire n297_o;
  wire n298_o;
  wire n299_o;
  wire n300_o;
  wire n301_o;
  wire [7:0] n306_o;
  wire [7:0] n307_o;
  wire [7:0] n308_o;
  wire [7:0] n309_o;
  wire [7:0] n310_o;
  wire [7:0] n311_o;
  wire [7:0] n312_o;
  wire [7:0] n313_o;
  wire [7:0] n314_o;
  wire [7:0] n315_o;
  wire [7:0] n316_o;
  wire [15:0] n317_o;
  wire [15:0] n318_o;
  wire [15:0] n319_o;
  wire [15:0] n320_o;
  wire [15:0] n321_o;
  wire [15:0] n322_o;
  wire [15:0] n323_o;
  wire [15:0] n324_o;
  wire [15:0] n325_o;
  wire [7:0] n326_o;
  wire [7:0] n327_o;
  wire [7:0] n328_o;
  wire [7:0] n329_o;
  wire [7:0] n330_o;
  wire [7:0] n331_o;
  wire [7:0] n332_o;
  wire [7:0] n333_o;
  wire [7:0] n334_o;
  wire n335_o;
  wire [15:0] n336_o;
  wire [15:0] n337_o;
  wire n338_o;
  wire n339_o;
  wire n340_o;
  wire n341_o;
  wire n342_o;
  wire n343_o;
  wire n345_o;
  wire n346_o;
  wire n349_o;
  wire n351_o;
  wire [1:0] n352_o;
  reg n355_o;
  reg n358_o;
  wire n361_o;
  wire n363_o;
  wire n365_o;
  wire n367_o;
  wire n369_o;
  wire n371_o;
  wire n373_o;
  wire n376_o;
  wire n379_o;
  wire n384_o;
  wire n385_o;
  wire [3:0] n386_o;
  wire n387_o;
  wire [2:0] n388_o;
  wire [3:0] n390_o;
  wire [2:0] n391_o;
  wire [3:0] n392_o;
  wire [3:0] n393_o;
  wire [2:0] n394_o;
  wire [3:0] n396_o;
  wire [2:0] n397_o;
  wire [3:0] n399_o;
  wire [2:0] n400_o;
  wire [3:0] n401_o;
  wire [2:0] n402_o;
  wire n404_o;
  wire n405_o;
  wire [2:0] n406_o;
  wire [3:0] n407_o;
  wire [2:0] n408_o;
  wire [3:0] n410_o;
  wire [3:0] n411_o;
  wire [3:0] n412_o;
  wire [3:0] n414_o;
  wire [3:0] n415_o;
  wire [3:0] n416_o;
  wire [3:0] n417_o;
  wire [3:0] n418_o;
  wire [3:0] n419_o;
  wire [3:0] n420_o;
  wire [3:0] n421_o;
  wire n425_o;
  wire n426_o;
  wire n427_o;
  wire [3:0] n429_o;
  wire [3:0] n430_o;
  wire [2:0] n431_o;
  wire [3:0] n433_o;
  wire [2:0] n434_o;
  wire [3:0] n436_o;
  wire [2:0] n437_o;
  wire [3:0] n439_o;
  wire [2:0] n440_o;
  wire [3:0] n442_o;
  wire [2:0] n443_o;
  wire [3:0] n445_o;
  wire [2:0] n446_o;
  wire [3:0] n447_o;
  wire n448_o;
  wire [2:0] n449_o;
  wire [3:0] n450_o;
  wire [3:0] n452_o;
  wire [3:0] n453_o;
  wire [3:0] n454_o;
  wire [3:0] n455_o;
  wire [3:0] n456_o;
  wire [3:0] n457_o;
  wire [3:0] n458_o;
  wire [3:0] n459_o;
  wire n463_o;
  wire n464_o;
  wire n465_o;
  wire n466_o;
  wire n467_o;
  wire n468_o;
  wire n469_o;
  wire n470_o;
  wire n471_o;
  wire [31:0] n472_o;
  wire [31:0] n473_o;
  wire [31:0] n475_o;
  wire [15:0] n479_o;
  wire n480_o;
  wire n481_o;
  wire n482_o;
  wire n483_o;
  wire n484_o;
  wire n485_o;
  wire n486_o;
  wire n487_o;
  wire n488_o;
  wire n489_o;
  wire n490_o;
  wire n491_o;
  wire n492_o;
  wire n493_o;
  wire n494_o;
  wire n495_o;
  wire [3:0] n496_o;
  wire [3:0] n497_o;
  wire [3:0] n498_o;
  wire [3:0] n499_o;
  wire [15:0] n500_o;
  wire n501_o;
  localparam [15:0] n502_o = 16'b1111111111111111;
  wire n503_o;
  wire n504_o;
  wire n505_o;
  wire n506_o;
  wire n507_o;
  wire n508_o;
  wire n509_o;
  wire n510_o;
  wire n511_o;
  wire n512_o;
  wire n513_o;
  wire [7:0] n514_o;
  wire n515_o;
  wire n516_o;
  wire n517_o;
  wire n518_o;
  wire n519_o;
  wire n520_o;
  wire n521_o;
  wire n522_o;
  wire [3:0] n523_o;
  wire [3:0] n524_o;
  wire [7:0] n525_o;
  wire n526_o;
  wire [2:0] n527_o;
  wire [2:0] n528_o;
  wire n530_o;
  wire n533_o;
  wire n536_o;
  wire n537_o;
  wire n538_o;
  wire n539_o;
  wire [15:0] n540_o;
  wire [15:0] n541_o;
  wire [15:0] n542_o;
  wire [15:0] n543_o;
  wire [15:0] n544_o;
  wire [31:0] n545_o;
  wire [15:0] n546_o;
  wire [15:0] n547_o;
  wire [15:0] n548_o;
  wire [15:0] n549_o;
  wire [15:0] n550_o;
  wire [31:0] n551_o;
  wire [31:0] n552_o;
  wire [31:0] n553_o;
  wire [15:0] n556_o;
  wire [15:0] n557_o;
  wire n558_o;
  wire n559_o;
  wire n560_o;
  wire n561_o;
  wire n562_o;
  wire n563_o;
  wire n564_o;
  wire n565_o;
  wire n566_o;
  wire n567_o;
  wire n568_o;
  wire n569_o;
  wire n570_o;
  wire n571_o;
  wire n572_o;
  wire n573_o;
  wire n574_o;
  wire n575_o;
  wire n576_o;
  wire n577_o;
  wire n578_o;
  wire n579_o;
  wire n580_o;
  wire n581_o;
  wire n582_o;
  wire [3:0] n583_o;
  wire [3:0] n584_o;
  wire [3:0] n585_o;
  wire [3:0] n586_o;
  wire [3:0] n587_o;
  wire [3:0] n588_o;
  wire [15:0] n589_o;
  wire [7:0] n590_o;
  wire [23:0] n591_o;
  wire [7:0] n592_o;
  wire [7:0] n593_o;
  wire [7:0] n594_o;
  wire [7:0] n595_o;
  wire [7:0] n596_o;
  wire [7:0] n597_o;
  wire [7:0] n598_o;
  wire [23:0] n599_o;
  wire [23:0] n600_o;
  wire [7:0] n601_o;
  wire [7:0] n602_o;
  wire [7:0] n603_o;
  wire [7:0] n604_o;
  wire [7:0] n605_o;
  wire [7:0] n606_o;
  wire [7:0] n607_o;
  wire n612_o;
  wire n614_o;
  wire n615_o;
  wire n616_o;
  wire n618_o;
  wire n620_o;
  wire n623_o;
  wire n625_o;
  wire n627_o;
  wire n628_o;
  wire n630_o;
  wire n631_o;
  wire n633_o;
  wire n635_o;
  wire n636_o;
  wire n637_o;
  wire n639_o;
  wire n641_o;
  wire n642_o;
  wire n644_o;
  wire n646_o;
  wire n648_o;
  wire n649_o;
  wire n651_o;
  wire n653_o;
  wire n654_o;
  wire n655_o;
  wire n656_o;
  wire n657_o;
  wire n658_o;
  wire n660_o;
  wire n661_o;
  wire n662_o;
  wire [31:0] n663_o;
  wire [31:0] n664_o;
  wire [31:0] n665_o;
  wire n666_o;
  wire n668_o;
  wire n669_o;
  wire n670_o;
  wire n671_o;
  wire n672_o;
  wire n674_o;
  wire [11:0] n675_o;
  wire [15:0] n677_o;
  wire [11:0] n678_o;
  wire [15:0] n680_o;
  wire n681_o;
  wire n682_o;
  wire n683_o;
  wire n684_o;
  wire [15:0] n685_o;
  wire n686_o;
  wire n687_o;
  wire n688_o;
  wire n689_o;
  wire n690_o;
  wire n692_o;
  wire n693_o;
  wire n694_o;
  wire [23:0] n695_o;
  wire [23:0] n696_o;
  wire [23:0] n697_o;
  wire [7:0] n698_o;
  wire n699_o;
  wire [15:0] n700_o;
  wire [15:0] n701_o;
  wire [15:0] n702_o;
  wire [15:0] n703_o;
  wire [15:0] n704_o;
  wire [15:0] n705_o;
  wire [15:0] n706_o;
  wire [31:0] n707_o;
  wire [31:0] n708_o;
  wire [15:0] n709_o;
  wire [15:0] n710_o;
  wire [15:0] n711_o;
  wire [15:0] n712_o;
  wire [15:0] n713_o;
  wire [31:0] n714_o;
  wire [31:0] n715_o;
  wire [31:0] n716_o;
  wire [31:0] n717_o;
  wire [31:0] n718_o;
  wire [31:0] n719_o;
  wire [31:0] n720_o;
  wire [15:0] n721_o;
  wire [15:0] n722_o;
  wire [15:0] n723_o;
  wire [15:0] n724_o;
  wire [15:0] n725_o;
  wire n726_o;
  wire [31:0] n727_o;
  wire [31:0] n728_o;
  wire n729_o;
  wire n732_o;
  wire [31:0] n733_o;
  wire n734_o;
  wire n736_o;
  wire [31:0] n737_o;
  wire n738_o;
  wire n740_o;
  wire [31:0] n742_o;
  wire [31:0] n743_o;
  wire n744_o;
  wire n745_o;
  wire n746_o;
  wire n747_o;
  wire n748_o;
  wire n749_o;
  wire n750_o;
  wire [31:0] n751_o;
  wire [31:0] n752_o;
  wire n754_o;
  wire n756_o;
  wire n757_o;
  wire n759_o;
  wire n761_o;
  wire n762_o;
  wire n764_o;
  wire n777_o;
  wire [15:0] n778_o;
  wire n779_o;
  wire n780_o;
  wire n781_o;
  wire n782_o;
  wire n783_o;
  wire n784_o;
  wire n785_o;
  wire n786_o;
  wire n787_o;
  wire n788_o;
  wire n789_o;
  wire n790_o;
  wire n791_o;
  wire n792_o;
  wire n793_o;
  wire n794_o;
  wire [3:0] n795_o;
  wire [3:0] n796_o;
  wire [3:0] n797_o;
  wire [3:0] n798_o;
  wire [15:0] n799_o;
  wire [15:0] n800_o;
  wire [15:0] n801_o;
  wire [31:0] n802_o;
  wire n803_o;
  wire n805_o;
  wire n807_o;
  wire [1:0] n808_o;
  wire [15:0] n809_o;
  wire [31:0] n810_o;
  wire n812_o;
  wire [14:0] n813_o;
  wire [15:0] n814_o;
  wire [30:0] n815_o;
  wire [31:0] n817_o;
  wire n819_o;
  wire [13:0] n820_o;
  wire [15:0] n821_o;
  wire [29:0] n822_o;
  wire [31:0] n824_o;
  wire n826_o;
  wire [12:0] n827_o;
  wire [15:0] n828_o;
  wire [28:0] n829_o;
  wire [31:0] n831_o;
  wire n833_o;
  wire [3:0] n834_o;
  reg [31:0] n835_o;
  wire [31:0] n836_o;
  wire [9:0] n843_o;
  wire [9:0] n844_o;
  wire [9:0] n846_o;
  wire [9:0] n848_o;
  wire [9:0] n850_o;
  wire n851_o;
  wire [9:0] n853_o;
  wire [9:0] n855_o;
  wire [9:0] n857_o;
  wire [9:0] n859_o;
  wire [9:0] n861_o;
  wire [9:0] n863_o;
  wire [3:0] n864_o;
  wire [7:0] n866_o;
  wire [9:0] n868_o;
  wire [9:0] n869_o;
  wire n870_o;
  wire [9:0] n872_o;
  wire [9:0] n873_o;
  wire [31:0] n874_o;
  wire [31:0] n877_o;
  wire [31:0] n878_o;
  wire n880_o;
  wire n881_o;
  wire n882_o;
  wire [2:0] n883_o;
  wire n884_o;
  wire n885_o;
  wire n886_o;
  wire n887_o;
  wire n888_o;
  wire n889_o;
  wire n890_o;
  wire n891_o;
  wire [3:0] n892_o;
  wire [3:0] n893_o;
  wire [7:0] n894_o;
  wire n895_o;
  wire n896_o;
  wire n897_o;
  wire n898_o;
  wire n899_o;
  wire n900_o;
  wire n901_o;
  wire n902_o;
  wire n903_o;
  wire n904_o;
  wire n905_o;
  wire n906_o;
  wire n907_o;
  wire n908_o;
  wire n909_o;
  wire n910_o;
  wire [3:0] n911_o;
  wire [3:0] n912_o;
  wire [3:0] n913_o;
  wire [3:0] n914_o;
  wire [15:0] n915_o;
  wire n916_o;
  wire [31:0] n917_o;
  wire [7:0] n918_o;
  wire [7:0] n919_o;
  wire [7:0] n920_o;
  wire [23:0] n921_o;
  wire [23:0] n922_o;
  wire [23:0] n923_o;
  wire [31:0] n924_o;
  wire [31:0] n925_o;
  wire n926_o;
  wire n927_o;
  wire n930_o;
  wire n931_o;
  wire n932_o;
  wire n933_o;
  wire [4:0] n936_o;
  wire [4:0] n937_o;
  wire [3:0] n939_o;
  wire [4:0] n941_o;
  wire [4:0] n942_o;
  wire [4:0] n943_o;
  wire [4:0] n944_o;
  wire [4:0] n945_o;
  wire [26:0] n946_o;
  wire [26:0] n947_o;
  wire [26:0] n948_o;
  wire n950_o;
  wire n952_o;
  wire n953_o;
  wire n954_o;
  wire n955_o;
  wire n957_o;
  wire n958_o;
  wire n959_o;
  wire n960_o;
  wire n961_o;
  wire n962_o;
  wire n963_o;
  wire n965_o;
  wire n966_o;
  wire n967_o;
  wire n969_o;
  wire n970_o;
  wire n971_o;
  wire n972_o;
  wire n973_o;
  wire n976_o;
  wire [31:0] n977_o;
  wire n979_o;
  wire [31:0] n980_o;
  wire [31:0] n982_o;
  wire n984_o;
  wire [31:0] n985_o;
  wire [31:0] n987_o;
  wire n989_o;
  wire [31:0] n990_o;
  wire [31:0] n992_o;
  wire n994_o;
  wire [31:0] n995_o;
  wire [31:0] n997_o;
  wire n999_o;
  wire [31:0] n1000_o;
  wire [31:0] n1002_o;
  wire n1004_o;
  wire [31:0] n1005_o;
  wire [31:0] n1007_o;
  wire n1009_o;
  wire [31:0] n1010_o;
  wire [31:0] n1012_o;
  wire n1015_o;
  wire n1017_o;
  wire n1018_o;
  wire n1019_o;
  wire n1020_o;
  wire n1021_o;
  wire n1023_o;
  wire n1024_o;
  wire [31:0] n1033_o;
  wire [31:0] n1034_o;
  wire [31:0] n1035_o;
  wire n1036_o;
  wire [31:0] n1038_o;
  wire [31:0] n1042_o;
  localparam [2:0] n1043_o = 3'b000;
  wire n1044_o;
  wire n1045_o;
  wire n1046_o;
  wire n1047_o;
  wire n1048_o;
  wire [3:0] n1049_o;
  wire n1050_o;
  wire n1051_o;
  wire n1052_o;
  wire n1053_o;
  wire n1054_o;
  wire n1055_o;
  wire n1056_o;
  wire n1057_o;
  wire [3:0] n1058_o;
  wire [3:0] n1059_o;
  wire [7:0] n1060_o;
  wire n1061_o;
  wire n1062_o;
  wire n1063_o;
  wire n1064_o;
  wire n1065_o;
  wire n1066_o;
  wire n1067_o;
  wire n1068_o;
  wire n1069_o;
  wire n1070_o;
  wire n1071_o;
  wire n1072_o;
  wire n1073_o;
  wire n1074_o;
  wire n1075_o;
  wire n1076_o;
  wire [3:0] n1077_o;
  wire [3:0] n1078_o;
  wire [3:0] n1079_o;
  wire [3:0] n1080_o;
  wire [15:0] n1081_o;
  localparam [1:0] n1082_o = 2'b11;
  wire n1085_o;
  wire n1086_o;
  wire n1090_o;
  wire n1091_o;
  wire n1092_o;
  wire n1093_o;
  wire n1094_o;
  wire n1095_o;
  wire n1096_o;
  wire n1097_o;
  wire n1098_o;
  wire n1099_o;
  wire n1100_o;
  wire n1101_o;
  wire n1102_o;
  wire n1103_o;
  wire n1104_o;
  wire n1105_o;
  wire n1107_o;
  wire n1109_o;
  wire n1111_o;
  wire n1112_o;
  wire n1113_o;
  wire n1114_o;
  wire [2:0] n1115_o;
  wire n1116_o;
  wire n1117_o;
  wire [1:0] n1118_o;
  wire n1119_o;
  wire n1120_o;
  wire n1121_o;
  wire [1:0] n1122_o;
  wire [1:0] n1123_o;
  wire [7:0] n1127_o;
  wire [7:0] n1128_o;
  wire [7:0] n1129_o;
  wire [23:0] n1130_o;
  wire [23:0] n1131_o;
  wire [23:0] n1132_o;
  wire [31:0] n1133_o;
  wire [31:0] n1134_o;
  wire [31:0] n1135_o;
  wire [31:0] n1136_o;
  wire n1138_o;
  wire n1140_o;
  wire n1141_o;
  wire n1142_o;
  wire n1143_o;
  wire n1144_o;
  wire n1146_o;
  wire n1147_o;
  wire n1148_o;
  wire n1150_o;
  wire n1151_o;
  wire n1152_o;
  wire n1153_o;
  wire n1154_o;
  wire [2:0] n1155_o;
  wire n1156_o;
  wire n1158_o;
  wire n1159_o;
  wire n1160_o;
  wire n1161_o;
  wire n1162_o;
  wire n1165_o;
  wire n1167_o;
  wire n1170_o;
  wire n1172_o;
  wire n1176_o;
  wire n1179_o;
  wire n1182_o;
  wire n1184_o;
  wire n1185_o;
  wire n1186_o;
  wire n1187_o;
  wire n1188_o;
  wire n1190_o;
  wire n1191_o;
  wire n1192_o;
  wire n1193_o;
  wire n1194_o;
  wire n1197_o;
  wire [2:0] n1199_o;
  wire [3:0] n1201_o;
  wire [5:0] n1203_o;
  wire [1:0] n1204_o;
  wire [1:0] n1205_o;
  wire [3:0] n1206_o;
  wire n1207_o;
  wire n1208_o;
  wire n1210_o;
  wire n1211_o;
  wire n1212_o;
  wire n1213_o;
  wire [31:0] n1214_o;
  wire [31:0] n1215_o;
  wire [31:0] n1216_o;
  wire [31:0] n1217_o;
  wire [5:0] n1218_o;
  wire [3:0] n1219_o;
  wire n1220_o;
  wire n1221_o;
  wire n1223_o;
  wire n1224_o;
  wire n1225_o;
  wire n1226_o;
  wire [7:0] n1228_o;
  wire n1231_o;
  wire n1234_o;
  wire [2:0] n1235_o;
  wire [7:0] n1236_o;
  wire n1238_o;
  wire n1242_o;
  wire n1245_o;
  wire [2:0] n1247_o;
  wire [7:0] n1248_o;
  wire n1249_o;
  wire n1250_o;
  wire n1251_o;
  wire n1253_o;
  wire [2:0] n1254_o;
  wire [7:0] n1255_o;
  wire n1257_o;
  wire n1258_o;
  wire n1259_o;
  wire [7:0] n1260_o;
  wire [7:0] n1261_o;
  wire n1263_o;
  wire [15:0] n1264_o;
  wire [31:0] n1265_o;
  wire [15:0] n1266_o;
  wire [7:0] n1267_o;
  wire n1269_o;
  wire [7:0] n1270_o;
  wire n1272_o;
  wire n1273_o;
  wire n1274_o;
  wire n1276_o;
  wire n1278_o;
  wire n1280_o;
  wire n1282_o;
  wire n1284_o;
  wire n1285_o;
  wire [31:0] n1286_o;
  wire [31:0] n1287_o;
  wire [31:0] n1289_o;
  wire [5:0] n1290_o;
  wire [5:0] n1291_o;
  wire [31:0] n1292_o;
  wire [5:0] n1293_o;
  wire n1294_o;
  wire n1295_o;
  wire n1296_o;
  wire n1297_o;
  wire n1298_o;
  wire n1299_o;
  wire n1300_o;
  wire n1301_o;
  wire n1302_o;
  wire n1303_o;
  wire n1304_o;
  wire [1:0] n1306_o;
  wire [1:0] n1307_o;
  wire n1309_o;
  wire n1311_o;
  wire n1312_o;
  wire n1313_o;
  wire n1314_o;
  wire n1316_o;
  wire n1318_o;
  wire n1320_o;
  wire n1321_o;
  wire n1322_o;
  wire n1323_o;
  wire n1325_o;
  wire n1326_o;
  wire n1328_o;
  wire n1329_o;
  wire n1330_o;
  wire n1331_o;
  wire n1332_o;
  wire n1333_o;
  wire n1334_o;
  wire n1335_o;
  wire n1338_o;
  wire n1339_o;
  wire n1340_o;
  wire n1342_o;
  wire n1343_o;
  wire n1344_o;
  wire n1345_o;
  wire n1348_o;
  wire [5:0] n1351_o;
  wire [5:0] n1354_o;
  wire n1356_o;
  wire [5:0] n1358_o;
  wire [5:0] n1360_o;
  wire n1362_o;
  wire [5:0] n1363_o;
  wire [5:0] n1364_o;
  wire n1365_o;
  wire [5:0] n1367_o;
  wire [5:0] n1369_o;
  wire n1370_o;
  wire [1:0] n1371_o;
  wire [1:0] n1373_o;
  wire n1375_o;
  wire [5:0] n1376_o;
  wire [5:0] n1377_o;
  wire n1378_o;
  wire [1:0] n1379_o;
  wire [1:0] n1381_o;
  wire n1383_o;
  wire [5:0] n1385_o;
  wire [5:0] n1386_o;
  wire n1387_o;
  wire n1388_o;
  wire n1390_o;
  wire [1:0] n1391_o;
  wire n1392_o;
  wire n1393_o;
  wire n1395_o;
  wire n1396_o;
  wire [5:0] n1397_o;
  wire n1398_o;
  wire n1399_o;
  wire n1400_o;
  wire n1401_o;
  wire n1403_o;
  wire n1405_o;
  wire n1406_o;
  wire [15:0] n1407_o;
  wire [15:0] n1408_o;
  wire [15:0] n1409_o;
  wire n1410_o;
  wire n1411_o;
  wire n1413_o;
  wire [15:0] n1414_o;
  wire [15:0] n1415_o;
  wire [31:0] n1416_o;
  wire n1417_o;
  wire n1418_o;
  wire n1420_o;
  wire [15:0] n1422_o;
  wire n1424_o;
  wire [15:0] n1425_o;
  wire [31:0] n1426_o;
  wire n1428_o;
  wire n1429_o;
  wire [7:0] n1430_o;
  wire [1:0] n1431_o;
  wire [1:0] n1432_o;
  wire [1:0] n1433_o;
  wire [1:0] n1434_o;
  wire n1435_o;
  wire [15:0] n1436_o;
  wire [15:0] n1437_o;
  wire n1438_o;
  wire n1439_o;
  wire n1440_o;
  wire n1441_o;
  wire n1442_o;
  wire n1443_o;
  wire n1444_o;
  wire n1445_o;
  wire n1446_o;
  wire n1447_o;
  wire n1448_o;
  wire n1449_o;
  wire n1450_o;
  wire n1451_o;
  wire n1452_o;
  wire n1453_o;
  wire n1454_o;
  wire n1455_o;
  wire n1456_o;
  wire n1457_o;
  wire [7:0] n1458_o;
  wire n1459_o;
  wire n1460_o;
  wire [5:0] n1461_o;
  wire [3:0] n1463_o;
  wire [5:0] n1464_o;
  wire n1465_o;
  wire n1466_o;
  wire n1467_o;
  wire n1468_o;
  wire n1469_o;
  wire [1:0] n1470_o;
  wire [1:0] n1471_o;
  wire [31:0] n1473_o;
  wire [1:0] n1475_o;
  wire [1:0] n1476_o;
  wire n1478_o;
  wire [15:0] n1480_o;
  wire [15:0] n1481_o;
  wire [31:0] n1482_o;
  wire [31:0] n1483_o;
  wire [15:0] n1485_o;
  wire n1486_o;
  wire n1488_o;
  wire [15:0] n1489_o;
  wire n1491_o;
  wire n1493_o;
  wire n1495_o;
  wire n1497_o;
  wire n1499_o;
  wire [1:0] n1500_o;
  wire [5:0] n1502_o;
  wire n1504_o;
  wire n1506_o;
  wire n1508_o;
  wire [7:0] n1509_o;
  wire n1511_o;
  wire n1513_o;
  wire [2:0] n1514_o;
  wire [7:0] n1515_o;
  wire n1517_o;
  wire n1519_o;
  wire [5:0] n1521_o;
  wire [3:0] n1522_o;
  wire [5:0] n1523_o;
  wire n1524_o;
  wire [5:0] n1525_o;
  wire [5:0] n1526_o;
  wire [31:0] n1527_o;
  wire [5:0] n1528_o;
  wire n1569_o;
  wire n1570_o;
  wire n1571_o;
  wire n1572_o;
  wire n1573_o;
  wire n1575_o;
  wire n1576_o;
  wire n1578_o;
  wire n1579_o;
  wire n1580_o;
  wire n1581_o;
  wire n1584_o;
  wire n1585_o;
  wire n1586_o;
  wire [1:0] n1587_o;
  wire n1588_o;
  wire n1589_o;
  wire n1590_o;
  wire [35:0] n1591_o;
  wire [47:0] n1592_o;
  wire [88:0] n1593_o;
  wire n1594_o;
  wire n1595_o;
  wire n1596_o;
  wire n1597_o;
  wire n1598_o;
  wire [84:0] n1600_o;
  wire n1601_o;
  wire n1602_o;
  wire n1603_o;
  wire n1604_o;
  wire n1605_o;
  wire [1:0] n1606_o;
  wire n1608_o;
  wire [88:0] n1610_o;
  wire [88:0] n1611_o;
  wire n1613_o;
  wire n1614_o;
  wire [16:0] n1615_o;
  wire [16:0] n1616_o;
  wire [16:0] n1617_o;
  wire [70:0] n1618_o;
  wire [70:0] n1619_o;
  wire [70:0] n1620_o;
  wire [88:0] n1622_o;
  wire n1630_o;
  wire [4:0] n1631_o;
  wire [5:0] n1633_o;
  wire [4:0] n1634_o;
  wire [5:0] n1636_o;
  wire n1638_o;
  wire [4:0] n1639_o;
  localparam [31:0] n1640_o = 32'b00000000000000000000000000000000;
  wire [26:0] n1641_o;
  wire [31:0] n1642_o;
  wire [31:0] n1643_o;
  wire n1645_o;
  wire [4:0] n1646_o;
  wire [4:0] n1648_o;
  wire [4:0] n1649_o;
  wire [4:0] n1651_o;
  wire [4:0] n1652_o;
  wire [5:0] n1653_o;
  wire n1654_o;
  wire n1655_o;
  wire [2:0] n1656_o;
  wire n1658_o;
  wire [5:0] n1660_o;
  wire [4:0] n1663_o;
  wire [4:0] n1664_o;
  wire [4:0] n1665_o;
  wire [1:0] n1666_o;
  wire n1668_o;
  wire [2:0] n1669_o;
  wire n1671_o;
  wire [5:0] n1673_o;
  wire [5:0] n1675_o;
  wire [4:0] n1678_o;
  wire [4:0] n1679_o;
  wire [4:0] n1680_o;
  wire [2:0] n1681_o;
  wire n1683_o;
  wire [2:0] n1684_o;
  wire [5:0] n1686_o;
  wire [5:0] n1688_o;
  wire [4:0] n1690_o;
  wire [2:0] n1691_o;
  wire [2:0] n1693_o;
  wire [5:0] n1695_o;
  wire [5:0] n1696_o;
  wire [5:0] n1697_o;
  wire [1:0] n1699_o;
  wire [1:0] n1700_o;
  wire [1:0] n1701_o;
  wire [1:0] n1702_o;
  wire n1703_o;
  wire n1704_o;
  wire n1705_o;
  wire [2:0] n1706_o;
  wire [2:0] n1707_o;
  wire [2:0] n1708_o;
  wire [5:0] n1709_o;
  wire [5:0] n1710_o;
  wire [2:0] n1711_o;
  wire n1713_o;
  wire n1715_o;
  wire n1717_o;
  wire n1719_o;
  wire [3:0] n1720_o;
  reg [5:0] n1726_o;
  wire n1728_o;
  wire [5:0] n1730_o;
  wire n1734_o;
  wire [7:0] n1735_o;
  wire [7:0] n1736_o;
  wire n1737_o;
  wire [7:0] n1738_o;
  wire [7:0] n1739_o;
  wire n1740_o;
  wire [7:0] n1741_o;
  wire [7:0] n1742_o;
  wire [7:0] n1743_o;
  wire [7:0] n1744_o;
  wire [7:0] n1745_o;
  wire [7:0] n1746_o;
  wire n1749_o;
  wire n1750_o;
  wire n1751_o;
  wire n1752_o;
  wire n1753_o;
  wire n1754_o;
  wire n1755_o;
  wire n1756_o;
  wire n1757_o;
  wire n1758_o;
  wire n1759_o;
  wire n1761_o;
  wire n1762_o;
  wire n1764_o;
  wire n1765_o;
  wire n1766_o;
  wire n1767_o;
  wire n1768_o;
  wire n1769_o;
  wire n1770_o;
  wire n1771_o;
  wire n1772_o;
  wire n1773_o;
  wire n1775_o;
  wire n1777_o;
  wire n1779_o;
  wire n1780_o;
  wire n1782_o;
  wire n1783_o;
  wire n1784_o;
  wire [4:0] n1786_o;
  wire n1787_o;
  wire [7:0] n1788_o;
  wire n1790_o;
  wire [2:0] n1791_o;
  wire [2:0] n1792_o;
  wire [2:0] n1793_o;
  wire [2:0] n1794_o;
  wire [4:0] n1795_o;
  wire [4:0] n1796_o;
  wire [4:0] n1797_o;
  wire n1798_o;
  wire n1799_o;
  wire n1800_o;
  wire n1801_o;
  wire n1802_o;
  wire n1803_o;
  wire [7:0] n1804_o;
  wire n1807_o;
  wire n1808_o;
  wire n1809_o;
  wire n1812_o;
  wire n1813_o;
  wire n1814_o;
  wire n1815_o;
  wire n1816_o;
  wire n1817_o;
  wire n1818_o;
  wire n1819_o;
  wire n1826_o;
  wire n1827_o;
  wire n1828_o;
  wire n1829_o;
  wire n1830_o;
  wire n1831_o;
  wire [2:0] n1833_o;
  wire [2:0] n1834_o;
  wire [2:0] n1835_o;
  wire n1836_o;
  wire n1837_o;
  wire [7:0] n1838_o;
  wire [7:0] n1839_o;
  wire n1840_o;
  wire n1841_o;
  wire n1842_o;
  wire n1843_o;
  wire [7:0] n1845_o;
  wire n1847_o;
  wire n1849_o;
  wire n1851_o;
  wire [1:0] n1861_o;
  wire n1863_o;
  wire [5:0] n1865_o;
  wire [5:0] n1867_o;
  localparam [88:0] n1870_o = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [1:0] n1873_o;
  wire n1875_o;
  wire n1877_o;
  wire [1:0] n1878_o;
  reg [1:0] n1882_o;
  wire n1883_o;
  wire n1885_o;
  wire n1886_o;
  wire n1889_o;
  wire n1890_o;
  wire n1892_o;
  wire n1893_o;
  wire [1:0] n1896_o;
  wire n1899_o;
  wire [6:0] n1904_o;
  wire n1906_o;
  wire n1907_o;
  wire n1908_o;
  wire n1909_o;
  wire n1910_o;
  wire n1911_o;
  wire n1912_o;
  wire [6:0] n1915_o;
  wire n1916_o;
  wire n1918_o;
  wire n1919_o;
  wire n1920_o;
  wire n1922_o;
  wire [1:0] n1924_o;
  wire n1926_o;
  wire n1927_o;
  wire [6:0] n1930_o;
  wire n1932_o;
  wire n1933_o;
  wire n1934_o;
  wire n1935_o;
  wire n1936_o;
  wire [6:0] n1939_o;
  wire n1940_o;
  wire n1942_o;
  wire [1:0] n1944_o;
  wire n1945_o;
  wire [6:0] n1946_o;
  wire n1948_o;
  wire n1949_o;
  wire n1950_o;
  wire n1951_o;
  wire n1953_o;
  wire [1:0] n1955_o;
  wire n1956_o;
  wire n1957_o;
  wire n1958_o;
  wire n1959_o;
  wire n1961_o;
  wire n1962_o;
  wire [1:0] n1965_o;
  wire n1966_o;
  wire [6:0] n1968_o;
  wire n1969_o;
  wire n1974_o;
  wire [1:0] n1976_o;
  wire [1:0] n1977_o;
  wire [1:0] n1978_o;
  wire n1981_o;
  wire n1982_o;
  wire n1983_o;
  wire [1:0] n1985_o;
  wire n1986_o;
  wire n1987_o;
  wire n1988_o;
  wire n1990_o;
  wire n1991_o;
  wire n1994_o;
  wire n1995_o;
  wire n1996_o;
  wire [2:0] n1997_o;
  wire n1999_o;
  wire [2:0] n2001_o;
  wire n2003_o;
  wire n2005_o;
  wire n2006_o;
  wire n2007_o;
  wire n2008_o;
  wire n2010_o;
  wire n2011_o;
  wire [2:0] n2013_o;
  wire n2015_o;
  wire n2017_o;
  wire n2018_o;
  wire n2019_o;
  wire n2020_o;
  wire n2022_o;
  wire n2024_o;
  wire n2025_o;
  wire n2027_o;
  wire n2028_o;
  wire n2030_o;
  wire n2032_o;
  wire [2:0] n2033_o;
  wire n2035_o;
  wire n2038_o;
  wire n2041_o;
  wire n2044_o;
  wire n2046_o;
  wire n2048_o;
  wire n2050_o;
  wire [4:0] n2051_o;
  reg n2054_o;
  reg n2057_o;
  reg n2060_o;
  reg n2064_o;
  reg n2068_o;
  wire n2069_o;
  reg n2070_o;
  reg n2071_o;
  reg [6:0] n2076_o;
  wire n2078_o;
  wire [3:0] n2079_o;
  reg n2082_o;
  reg n2085_o;
  reg n2087_o;
  reg n2089_o;
  reg n2091_o;
  wire n2092_o;
  reg n2093_o;
  wire n2094_o;
  reg n2095_o;
  wire n2096_o;
  reg n2097_o;
  wire n2098_o;
  reg n2099_o;
  wire n2100_o;
  reg n2101_o;
  reg n2102_o;
  reg [6:0] n2105_o;
  wire n2107_o;
  wire n2110_o;
  wire n2113_o;
  wire n2116_o;
  wire n2119_o;
  wire [1:0] n2121_o;
  wire n2122_o;
  wire n2123_o;
  wire [1:0] n2124_o;
  wire [1:0] n2125_o;
  wire n2126_o;
  wire n2127_o;
  wire n2128_o;
  wire n2129_o;
  wire n2130_o;
  wire [1:0] n2136_o;
  wire [1:0] n2137_o;
  wire [6:0] n2139_o;
  wire [3:0] n2140_o;
  wire n2141_o;
  wire [2:0] n2142_o;
  wire n2144_o;
  wire n2145_o;
  wire n2148_o;
  wire n2149_o;
  wire n2153_o;
  wire n2154_o;
  wire n2156_o;
  wire n2158_o;
  wire n2159_o;
  wire n2161_o;
  wire n2162_o;
  wire n2163_o;
  wire n2165_o;
  wire n2166_o;
  wire n2167_o;
  wire [6:0] n2169_o;
  wire n2172_o;
  wire n2173_o;
  wire [2:0] n2174_o;
  wire n2176_o;
  wire n2177_o;
  wire [2:0] n2178_o;
  wire n2180_o;
  wire [5:0] n2181_o;
  wire n2183_o;
  wire n2184_o;
  wire n2185_o;
  wire n2186_o;
  wire n2187_o;
  wire [6:0] n2188_o;
  wire n2190_o;
  wire [1:0] n2191_o;
  wire n2193_o;
  wire n2194_o;
  wire n2195_o;
  wire [1:0] n2196_o;
  wire n2198_o;
  wire [2:0] n2199_o;
  wire n2201_o;
  wire n2202_o;
  wire [1:0] n2203_o;
  wire n2205_o;
  wire n2206_o;
  wire n2207_o;
  wire [1:0] n2210_o;
  wire n2212_o;
  wire [1:0] n2213_o;
  wire n2215_o;
  wire n2218_o;
  wire n2221_o;
  wire n2223_o;
  wire [1:0] n2224_o;
  wire n2226_o;
  wire [1:0] n2229_o;
  wire n2230_o;
  wire n2231_o;
  wire n2234_o;
  wire n2235_o;
  wire n2236_o;
  wire n2237_o;
  wire [6:0] n2239_o;
  wire n2242_o;
  wire n2244_o;
  wire n2246_o;
  wire n2247_o;
  wire [1:0] n2248_o;
  wire n2250_o;
  wire n2253_o;
  wire n2256_o;
  wire n2258_o;
  wire n2260_o;
  wire n2262_o;
  wire n2264_o;
  wire n2266_o;
  wire n2268_o;
  wire n2269_o;
  wire [2:0] n2270_o;
  wire n2272_o;
  wire n2273_o;
  wire n2274_o;
  wire [1:0] n2275_o;
  wire n2277_o;
  wire [1:0] n2278_o;
  wire n2280_o;
  wire n2281_o;
  wire [2:0] n2282_o;
  wire n2284_o;
  wire [1:0] n2285_o;
  wire n2287_o;
  wire n2288_o;
  wire n2289_o;
  wire n2290_o;
  wire [5:0] n2291_o;
  wire n2293_o;
  wire n2294_o;
  wire n2295_o;
  wire [1:0] n2296_o;
  wire n2298_o;
  wire n2300_o;
  wire [1:0] n2301_o;
  reg [1:0] n2305_o;
  wire n2306_o;
  wire [5:0] n2307_o;
  wire n2309_o;
  wire n2310_o;
  wire n2312_o;
  wire n2313_o;
  wire [6:0] n2315_o;
  wire n2318_o;
  wire n2319_o;
  wire n2320_o;
  wire n2321_o;
  wire [6:0] n2323_o;
  wire n2325_o;
  wire n2326_o;
  wire [1:0] n2332_o;
  wire n2335_o;
  wire n2336_o;
  wire n2337_o;
  wire n2338_o;
  wire n2339_o;
  wire n2340_o;
  wire n2341_o;
  wire n2342_o;
  wire n2343_o;
  wire [6:0] n2345_o;
  wire [1:0] n2346_o;
  wire n2348_o;
  wire n2349_o;
  wire n2350_o;
  wire n2351_o;
  wire n2352_o;
  wire n2353_o;
  wire n2354_o;
  wire n2355_o;
  wire n2356_o;
  wire n2357_o;
  wire n2358_o;
  wire n2359_o;
  wire [6:0] n2360_o;
  wire [1:0] n2361_o;
  wire [1:0] n2362_o;
  wire n2364_o;
  wire n2367_o;
  wire n2370_o;
  wire n2371_o;
  wire n2372_o;
  wire n2373_o;
  wire n2374_o;
  wire n2375_o;
  wire n2376_o;
  wire n2377_o;
  wire n2378_o;
  wire n2379_o;
  wire n2380_o;
  wire n2381_o;
  wire n2382_o;
  wire [6:0] n2383_o;
  wire [1:0] n2384_o;
  wire n2386_o;
  wire [1:0] n2387_o;
  wire n2389_o;
  wire n2390_o;
  wire [2:0] n2391_o;
  wire n2393_o;
  wire n2394_o;
  wire [2:0] n2395_o;
  wire n2397_o;
  wire n2398_o;
  wire [3:0] n2399_o;
  wire n2401_o;
  wire n2402_o;
  wire [1:0] n2404_o;
  wire n2407_o;
  wire n2408_o;
  wire n2409_o;
  wire n2410_o;
  wire [6:0] n2412_o;
  wire n2413_o;
  wire n2416_o;
  wire n2417_o;
  wire n2418_o;
  wire n2419_o;
  wire n2421_o;
  wire n2422_o;
  wire n2425_o;
  wire n2428_o;
  wire [1:0] n2430_o;
  wire n2432_o;
  wire n2433_o;
  wire n2434_o;
  wire [6:0] n2436_o;
  wire [1:0] n2437_o;
  wire n2438_o;
  wire n2441_o;
  wire n2444_o;
  wire n2446_o;
  wire [1:0] n2447_o;
  wire n2449_o;
  wire [1:0] n2450_o;
  wire [1:0] n2451_o;
  wire n2453_o;
  wire n2455_o;
  wire n2457_o;
  wire [6:0] n2458_o;
  wire [1:0] n2459_o;
  wire [1:0] n2460_o;
  wire n2462_o;
  wire n2463_o;
  wire n2464_o;
  wire n2466_o;
  wire n2468_o;
  wire n2469_o;
  wire n2470_o;
  wire n2471_o;
  wire n2472_o;
  wire n2473_o;
  wire n2474_o;
  wire n2475_o;
  wire n2476_o;
  wire n2477_o;
  wire n2479_o;
  wire n2480_o;
  wire n2481_o;
  wire n2482_o;
  wire n2484_o;
  wire n2486_o;
  wire [6:0] n2487_o;
  wire [1:0] n2488_o;
  wire [1:0] n2489_o;
  wire n2491_o;
  wire n2493_o;
  wire n2495_o;
  wire n2497_o;
  wire [1:0] n2498_o;
  wire [1:0] n2499_o;
  wire n2501_o;
  wire n2502_o;
  wire n2503_o;
  wire [1:0] n2504_o;
  wire [1:0] n2505_o;
  wire [1:0] n2506_o;
  wire [1:0] n2507_o;
  wire n2508_o;
  wire n2509_o;
  wire n2510_o;
  wire n2511_o;
  wire n2513_o;
  wire n2515_o;
  wire [6:0] n2516_o;
  wire [2:0] n2517_o;
  wire n2519_o;
  wire n2520_o;
  wire [1:0] n2521_o;
  wire n2523_o;
  wire n2524_o;
  wire [1:0] n2525_o;
  wire n2527_o;
  wire n2528_o;
  wire [2:0] n2529_o;
  wire n2531_o;
  wire [1:0] n2532_o;
  wire n2534_o;
  wire n2535_o;
  wire n2536_o;
  wire n2539_o;
  wire n2542_o;
  wire n2544_o;
  wire n2546_o;
  wire [1:0] n2547_o;
  wire n2549_o;
  wire [2:0] n2550_o;
  wire n2552_o;
  wire n2553_o;
  wire [2:0] n2554_o;
  wire n2556_o;
  wire [2:0] n2557_o;
  wire n2559_o;
  wire [1:0] n2560_o;
  wire n2562_o;
  wire n2563_o;
  wire [2:0] n2564_o;
  wire n2566_o;
  wire n2567_o;
  wire n2568_o;
  wire n2569_o;
  wire n2570_o;
  wire n2574_o;
  wire n2577_o;
  wire n2579_o;
  wire n2581_o;
  wire n2583_o;
  wire n2585_o;
  wire [2:0] n2586_o;
  wire n2588_o;
  wire [2:0] n2589_o;
  wire n2591_o;
  wire [1:0] n2592_o;
  wire n2594_o;
  wire n2595_o;
  wire [2:0] n2596_o;
  wire n2598_o;
  wire n2599_o;
  wire n2600_o;
  wire n2601_o;
  wire n2602_o;
  wire n2605_o;
  wire n2607_o;
  wire n2609_o;
  wire n2610_o;
  wire n2611_o;
  wire n2613_o;
  wire [2:0] n2614_o;
  wire n2616_o;
  wire [2:0] n2617_o;
  wire n2619_o;
  wire n2620_o;
  wire [2:0] n2621_o;
  wire n2623_o;
  wire [1:0] n2624_o;
  wire n2626_o;
  wire n2627_o;
  wire n2630_o;
  wire n2632_o;
  wire n2634_o;
  wire n2635_o;
  wire n2636_o;
  wire n2638_o;
  wire [2:0] n2639_o;
  wire n2641_o;
  wire [2:0] n2642_o;
  wire n2644_o;
  wire [1:0] n2645_o;
  wire n2647_o;
  wire n2648_o;
  wire [2:0] n2649_o;
  wire n2651_o;
  wire n2652_o;
  wire n2653_o;
  wire n2654_o;
  wire n2655_o;
  wire n2658_o;
  wire n2660_o;
  wire n2662_o;
  wire n2663_o;
  wire n2664_o;
  wire n2666_o;
  wire [2:0] n2667_o;
  wire n2669_o;
  wire [2:0] n2670_o;
  wire n2672_o;
  wire n2673_o;
  wire n2674_o;
  wire n2675_o;
  wire n2678_o;
  wire n2680_o;
  wire n2682_o;
  wire n2683_o;
  wire n2684_o;
  wire n2686_o;
  wire n2687_o;
  wire n2688_o;
  wire n2689_o;
  wire n2690_o;
  wire n2691_o;
  wire n2692_o;
  wire n2693_o;
  wire n2694_o;
  wire n2695_o;
  wire n2696_o;
  wire n2697_o;
  wire [5:0] n2698_o;
  wire n2700_o;
  wire n2701_o;
  wire n2702_o;
  wire n2703_o;
  wire n2704_o;
  wire n2705_o;
  wire n2706_o;
  wire n2707_o;
  wire n2708_o;
  wire n2709_o;
  wire n2710_o;
  wire n2711_o;
  wire n2713_o;
  wire n2715_o;
  wire n2716_o;
  wire n2718_o;
  wire n2719_o;
  wire n2720_o;
  wire [1:0] n2722_o;
  wire [2:0] n2723_o;
  wire [1:0] n2724_o;
  wire [2:0] n2725_o;
  wire [2:0] n2726_o;
  wire [1:0] n2727_o;
  wire [1:0] n2728_o;
  wire [6:0] n2730_o;
  wire [1:0] n2731_o;
  wire n2734_o;
  wire n2736_o;
  wire [2:0] n2737_o;
  wire [2:0] n2738_o;
  wire n2739_o;
  wire n2740_o;
  wire [1:0] n2741_o;
  wire [1:0] n2742_o;
  wire [6:0] n2743_o;
  wire n2744_o;
  wire n2745_o;
  wire [5:0] n2746_o;
  wire n2748_o;
  wire n2749_o;
  wire n2750_o;
  wire n2751_o;
  wire n2752_o;
  wire n2753_o;
  wire n2754_o;
  wire n2755_o;
  wire n2756_o;
  wire n2760_o;
  wire n2762_o;
  wire n2764_o;
  wire n2765_o;
  wire n2766_o;
  wire n2767_o;
  wire n2768_o;
  wire n2769_o;
  wire [6:0] n2771_o;
  wire [1:0] n2772_o;
  wire n2774_o;
  wire n2777_o;
  wire [2:0] n2778_o;
  wire n2780_o;
  wire [1:0] n2781_o;
  wire n2783_o;
  wire n2786_o;
  wire n2789_o;
  wire n2791_o;
  wire [1:0] n2792_o;
  wire n2794_o;
  wire n2796_o;
  wire n2797_o;
  wire n2799_o;
  wire n2800_o;
  wire n2802_o;
  wire n2804_o;
  wire n2806_o;
  wire n2808_o;
  wire n2810_o;
  wire n2811_o;
  wire n2813_o;
  wire n2815_o;
  wire n2816_o;
  wire [1:0] n2817_o;
  wire n2819_o;
  wire n2820_o;
  wire n2821_o;
  wire n2823_o;
  wire n2824_o;
  wire [2:0] n2825_o;
  wire [2:0] n2826_o;
  wire n2827_o;
  wire n2828_o;
  wire n2829_o;
  wire n2830_o;
  wire [1:0] n2831_o;
  wire [1:0] n2832_o;
  wire n2833_o;
  wire n2834_o;
  wire n2835_o;
  wire n2836_o;
  wire n2837_o;
  wire n2839_o;
  wire n2841_o;
  wire [6:0] n2842_o;
  wire n2843_o;
  wire n2845_o;
  wire n2846_o;
  wire n2848_o;
  wire n2850_o;
  wire n2852_o;
  wire n2854_o;
  wire n2855_o;
  wire n2856_o;
  wire n2858_o;
  wire n2860_o;
  wire n2861_o;
  wire n2862_o;
  wire n2863_o;
  wire n2864_o;
  wire n2865_o;
  wire n2867_o;
  wire n2869_o;
  wire [6:0] n2870_o;
  wire n2871_o;
  wire n2873_o;
  wire n2874_o;
  wire n2876_o;
  wire n2878_o;
  wire n2880_o;
  wire n2882_o;
  wire n2884_o;
  wire n2886_o;
  wire n2888_o;
  wire n2890_o;
  wire n2892_o;
  wire n2893_o;
  wire [3:0] n2894_o;
  wire n2896_o;
  wire [3:0] n2898_o;
  wire n2900_o;
  wire n2902_o;
  wire n2903_o;
  wire [1:0] n2904_o;
  wire n2906_o;
  wire n2907_o;
  wire n2908_o;
  wire n2909_o;
  wire n2911_o;
  wire [2:0] n2912_o;
  wire [2:0] n2913_o;
  wire n2914_o;
  wire n2915_o;
  wire n2916_o;
  wire n2917_o;
  wire [1:0] n2918_o;
  wire [1:0] n2919_o;
  wire n2920_o;
  wire n2921_o;
  wire n2922_o;
  wire n2923_o;
  wire n2924_o;
  wire n2926_o;
  wire [3:0] n2928_o;
  wire n2930_o;
  wire n2932_o;
  wire [6:0] n2933_o;
  wire n2934_o;
  wire [1:0] n2935_o;
  wire n2937_o;
  wire n2939_o;
  wire n2940_o;
  wire n2941_o;
  wire n2943_o;
  wire n2944_o;
  wire n2946_o;
  wire [2:0] n2947_o;
  wire [2:0] n2948_o;
  wire n2950_o;
  wire n2952_o;
  wire n2953_o;
  wire n2954_o;
  wire n2955_o;
  wire n2956_o;
  wire n2957_o;
  wire n2958_o;
  wire n2959_o;
  wire [1:0] n2960_o;
  wire [1:0] n2961_o;
  wire n2962_o;
  wire n2963_o;
  wire n2964_o;
  wire n2965_o;
  wire n2966_o;
  wire n2967_o;
  wire n2968_o;
  wire n2970_o;
  wire n2972_o;
  wire n2974_o;
  wire n2976_o;
  wire [3:0] n2978_o;
  wire n2980_o;
  wire n2982_o;
  wire [6:0] n2983_o;
  wire [1:0] n2984_o;
  wire [1:0] n2985_o;
  wire n2986_o;
  wire n2988_o;
  wire n2989_o;
  wire n2990_o;
  wire n2992_o;
  wire n2993_o;
  wire n2995_o;
  wire n2997_o;
  wire [1:0] n2998_o;
  wire [1:0] n2999_o;
  wire [2:0] n3000_o;
  wire [2:0] n3001_o;
  wire n3002_o;
  wire n3003_o;
  wire n3004_o;
  wire n3005_o;
  wire n3006_o;
  wire n3007_o;
  wire n3008_o;
  wire n3009_o;
  wire n3010_o;
  wire n3011_o;
  wire n3012_o;
  wire [1:0] n3013_o;
  wire [1:0] n3014_o;
  wire [1:0] n3015_o;
  wire [1:0] n3016_o;
  wire n3017_o;
  wire n3018_o;
  wire n3019_o;
  wire n3020_o;
  wire n3021_o;
  wire n3022_o;
  wire n3023_o;
  wire n3024_o;
  wire n3026_o;
  wire [3:0] n3028_o;
  wire n3030_o;
  wire n3031_o;
  wire n3032_o;
  wire [6:0] n3033_o;
  wire [1:0] n3035_o;
  wire [1:0] n3036_o;
  wire n3038_o;
  wire n3040_o;
  wire n3042_o;
  wire n3043_o;
  wire n3045_o;
  wire n3047_o;
  wire n3049_o;
  wire n3051_o;
  wire n3053_o;
  wire [1:0] n3054_o;
  wire [1:0] n3055_o;
  wire [2:0] n3056_o;
  wire [2:0] n3057_o;
  wire n3058_o;
  wire n3059_o;
  wire n3060_o;
  wire n3061_o;
  wire n3062_o;
  wire n3063_o;
  wire [1:0] n3064_o;
  wire [1:0] n3065_o;
  wire n3066_o;
  wire n3067_o;
  wire n3068_o;
  wire n3069_o;
  wire [1:0] n3070_o;
  wire [1:0] n3071_o;
  wire [1:0] n3072_o;
  wire [1:0] n3073_o;
  wire n3074_o;
  wire n3075_o;
  wire n3076_o;
  wire n3077_o;
  wire n3078_o;
  wire n3079_o;
  wire n3080_o;
  wire n3081_o;
  wire n3082_o;
  wire n3084_o;
  wire n3086_o;
  wire [3:0] n3088_o;
  wire n3090_o;
  wire n3092_o;
  wire n3093_o;
  wire [6:0] n3094_o;
  wire n3096_o;
  wire [1:0] n3097_o;
  wire n3099_o;
  wire [2:0] n3100_o;
  wire n3102_o;
  wire n3103_o;
  wire [3:0] n3104_o;
  wire n3106_o;
  wire [1:0] n3107_o;
  wire n3109_o;
  wire n3110_o;
  wire n3111_o;
  wire n3112_o;
  wire [2:0] n3113_o;
  wire n3115_o;
  wire [2:0] n3116_o;
  wire n3118_o;
  wire n3119_o;
  wire n3120_o;
  wire n3121_o;
  wire [2:0] n3123_o;
  wire n3125_o;
  wire n3127_o;
  wire n3128_o;
  wire [1:0] n3129_o;
  wire n3131_o;
  wire [1:0] n3132_o;
  wire n3134_o;
  wire n3137_o;
  wire n3139_o;
  wire [1:0] n3140_o;
  wire n3142_o;
  wire n3144_o;
  wire [1:0] n3145_o;
  reg [1:0] n3149_o;
  wire n3150_o;
  wire n3153_o;
  wire [1:0] n3154_o;
  wire n3156_o;
  wire n3157_o;
  wire [2:0] n3158_o;
  wire n3160_o;
  wire n3163_o;
  wire n3165_o;
  wire n3168_o;
  wire n3170_o;
  wire [1:0] n3171_o;
  wire n3173_o;
  wire n3174_o;
  wire n3175_o;
  wire n3176_o;
  wire [2:0] n3177_o;
  wire n3180_o;
  wire n3182_o;
  wire n3183_o;
  wire n3184_o;
  wire [2:0] n3186_o;
  wire n3188_o;
  wire n3190_o;
  wire n3191_o;
  wire n3192_o;
  wire n3193_o;
  wire n3194_o;
  wire n3195_o;
  wire n3196_o;
  wire [2:0] n3198_o;
  wire n3200_o;
  wire n3202_o;
  wire n3203_o;
  wire n3204_o;
  wire n3205_o;
  wire n3206_o;
  wire n3207_o;
  wire n3208_o;
  wire n3210_o;
  wire n3211_o;
  wire n3213_o;
  wire n3215_o;
  wire n3216_o;
  wire n3218_o;
  wire n3219_o;
  wire n3221_o;
  wire n3223_o;
  wire [2:0] n3224_o;
  wire n3226_o;
  wire n3229_o;
  wire [1:0] n3230_o;
  reg n3231_o;
  reg [6:0] n3234_o;
  wire n3236_o;
  wire [4:0] n3237_o;
  reg [1:0] n3239_o;
  reg n3241_o;
  wire n3242_o;
  reg n3243_o;
  wire n3244_o;
  wire n3245_o;
  wire n3246_o;
  reg n3247_o;
  wire n3248_o;
  wire n3249_o;
  wire n3250_o;
  reg n3251_o;
  reg n3252_o;
  reg n3253_o;
  reg n3254_o;
  reg [6:0] n3258_o;
  wire [1:0] n3259_o;
  wire n3260_o;
  wire [1:0] n3261_o;
  wire n3262_o;
  wire n3263_o;
  wire [1:0] n3264_o;
  wire n3265_o;
  wire n3266_o;
  wire n3267_o;
  wire [6:0] n3268_o;
  wire [1:0] n3269_o;
  wire n3270_o;
  wire n3271_o;
  wire n3273_o;
  wire n3276_o;
  wire n3278_o;
  wire n3280_o;
  wire n3283_o;
  wire n3286_o;
  wire n3289_o;
  wire [1:0] n3290_o;
  wire n3292_o;
  wire n3293_o;
  wire n3294_o;
  wire [1:0] n3295_o;
  wire [1:0] n3296_o;
  wire n3297_o;
  wire n3299_o;
  wire n3301_o;
  wire n3302_o;
  wire n3304_o;
  wire n3306_o;
  wire n3307_o;
  wire n3309_o;
  wire n3310_o;
  wire n3311_o;
  wire n3312_o;
  wire [2:0] n3313_o;
  wire n3315_o;
  wire [2:0] n3316_o;
  wire n3318_o;
  wire n3319_o;
  wire n3320_o;
  wire n3321_o;
  wire n3322_o;
  wire n3329_o;
  wire n3332_o;
  wire n3335_o;
  wire n3337_o;
  wire n3339_o;
  wire n3341_o;
  wire n3343_o;
  wire n3344_o;
  wire n3345_o;
  wire [1:0] n3346_o;
  wire n3348_o;
  wire n3349_o;
  wire n3350_o;
  wire [2:0] n3351_o;
  wire n3353_o;
  wire n3354_o;
  wire [3:0] n3355_o;
  wire n3357_o;
  wire n3358_o;
  wire [2:0] n3362_o;
  wire n3364_o;
  wire n3367_o;
  wire n3370_o;
  wire n3373_o;
  wire n3374_o;
  wire [1:0] n3376_o;
  wire n3378_o;
  wire n3380_o;
  wire n3382_o;
  wire n3383_o;
  wire n3386_o;
  wire n3389_o;
  wire n3392_o;
  wire n3394_o;
  wire n3396_o;
  wire n3397_o;
  wire n3400_o;
  wire n3403_o;
  wire n3405_o;
  wire n3406_o;
  wire n3407_o;
  wire n3409_o;
  wire n3411_o;
  wire [1:0] n3412_o;
  wire n3414_o;
  wire n3416_o;
  wire n3417_o;
  wire n3419_o;
  wire n3421_o;
  wire n3422_o;
  wire n3423_o;
  wire n3424_o;
  wire n3426_o;
  wire n3427_o;
  wire n3428_o;
  wire n3429_o;
  wire n3431_o;
  wire n3432_o;
  wire n3434_o;
  wire [2:0] n3435_o;
  wire n3437_o;
  wire [3:0] n3438_o;
  wire n3440_o;
  wire [1:0] n3441_o;
  wire n3443_o;
  wire n3444_o;
  wire n3445_o;
  wire n3446_o;
  wire n3448_o;
  wire n3449_o;
  wire n3450_o;
  wire n3451_o;
  wire n3452_o;
  wire n3453_o;
  wire n3454_o;
  wire n3455_o;
  wire n3458_o;
  wire n3459_o;
  wire n3461_o;
  wire n3462_o;
  wire n3463_o;
  wire n3464_o;
  wire n3465_o;
  wire n3466_o;
  wire n3467_o;
  wire n3468_o;
  wire n3471_o;
  wire [1:0] n3473_o;
  wire n3476_o;
  wire n3478_o;
  wire n3479_o;
  wire n3480_o;
  wire [1:0] n3482_o;
  wire n3484_o;
  wire n3485_o;
  wire n3486_o;
  wire n3487_o;
  wire n3488_o;
  wire n3489_o;
  wire [1:0] n3490_o;
  wire n3492_o;
  wire n3493_o;
  wire n3494_o;
  wire n3495_o;
  wire n3496_o;
  wire n3498_o;
  wire n3499_o;
  wire n3502_o;
  wire n3506_o;
  wire n3509_o;
  wire n3511_o;
  wire n3513_o;
  wire n3516_o;
  wire n3517_o;
  wire n3518_o;
  wire n3520_o;
  wire [1:0] n3521_o;
  wire n3523_o;
  wire n3525_o;
  wire n3527_o;
  wire n3529_o;
  wire n3531_o;
  wire n3532_o;
  wire n3533_o;
  wire n3535_o;
  wire n3537_o;
  wire [1:0] n3538_o;
  wire [1:0] n3539_o;
  wire n3541_o;
  wire n3543_o;
  wire n3544_o;
  wire n3546_o;
  wire n3547_o;
  wire n3548_o;
  wire n3549_o;
  wire n3550_o;
  wire n3551_o;
  wire n3552_o;
  wire n3553_o;
  wire n3554_o;
  wire n3555_o;
  wire n3556_o;
  wire n3557_o;
  wire n3559_o;
  wire n3561_o;
  wire n3563_o;
  wire n3565_o;
  wire n3567_o;
  wire [2:0] n3568_o;
  wire [2:0] n3569_o;
  wire n3571_o;
  wire [2:0] n3572_o;
  wire n3574_o;
  wire [1:0] n3575_o;
  wire n3577_o;
  wire n3578_o;
  wire n3579_o;
  wire [1:0] n3580_o;
  wire n3582_o;
  wire n3583_o;
  wire n3584_o;
  wire n3586_o;
  wire n3588_o;
  wire n3589_o;
  wire n3591_o;
  wire n3593_o;
  wire n3594_o;
  wire n3595_o;
  wire n3596_o;
  wire n3598_o;
  wire [1:0] n3599_o;
  wire n3601_o;
  wire n3604_o;
  wire n3605_o;
  wire [1:0] n3607_o;
  wire n3610_o;
  wire n3613_o;
  wire n3616_o;
  wire n3619_o;
  wire n3621_o;
  wire n3623_o;
  wire [1:0] n3627_o;
  wire n3629_o;
  wire n3632_o;
  wire n3634_o;
  wire n3635_o;
  wire n3636_o;
  wire n3637_o;
  wire n3639_o;
  wire n3642_o;
  wire n3644_o;
  wire n3646_o;
  wire n3648_o;
  wire n3649_o;
  wire n3650_o;
  wire n3651_o;
  wire n3652_o;
  wire n3654_o;
  wire n3656_o;
  wire n3658_o;
  wire n3659_o;
  wire n3660_o;
  wire n3661_o;
  wire n3663_o;
  wire n3665_o;
  wire n3668_o;
  wire n3670_o;
  wire n3672_o;
  wire n3674_o;
  wire n3675_o;
  wire n3676_o;
  wire n3677_o;
  wire n3678_o;
  wire [1:0] n3679_o;
  wire [1:0] n3681_o;
  wire n3683_o;
  wire n3685_o;
  wire n3687_o;
  wire [2:0] n3688_o;
  wire n3690_o;
  wire [2:0] n3691_o;
  wire n3693_o;
  wire [1:0] n3694_o;
  wire n3696_o;
  wire n3697_o;
  wire n3698_o;
  wire [1:0] n3699_o;
  wire n3701_o;
  wire n3702_o;
  wire n3704_o;
  wire n3706_o;
  wire [1:0] n3708_o;
  wire n3710_o;
  wire n3713_o;
  wire [1:0] n3715_o;
  wire n3718_o;
  wire n3721_o;
  wire n3724_o;
  wire n3727_o;
  wire n3729_o;
  wire n3731_o;
  wire n3733_o;
  wire n3735_o;
  wire n3736_o;
  wire n3737_o;
  wire n3738_o;
  wire n3740_o;
  wire n3742_o;
  wire n3743_o;
  wire [1:0] n3744_o;
  wire n3746_o;
  wire n3749_o;
  wire n3750_o;
  wire n3751_o;
  wire n3753_o;
  wire n3755_o;
  wire n3757_o;
  wire n3759_o;
  wire n3760_o;
  wire n3761_o;
  wire n3763_o;
  wire n3765_o;
  wire n3766_o;
  wire n3767_o;
  wire n3768_o;
  wire n3770_o;
  wire n3772_o;
  wire n3774_o;
  wire n3776_o;
  wire n3777_o;
  wire n3778_o;
  wire n3780_o;
  wire n3782_o;
  wire n3784_o;
  wire n3786_o;
  wire [1:0] n3787_o;
  wire n3789_o;
  wire [2:0] n3790_o;
  wire n3792_o;
  wire [3:0] n3793_o;
  wire n3795_o;
  wire [1:0] n3796_o;
  wire n3798_o;
  wire n3799_o;
  wire n3800_o;
  wire [1:0] n3801_o;
  wire n3803_o;
  wire n3804_o;
  wire n3806_o;
  wire n3807_o;
  wire n3808_o;
  wire n3809_o;
  wire n3810_o;
  wire n3812_o;
  wire n3813_o;
  wire [1:0] n3815_o;
  wire n3818_o;
  wire n3821_o;
  wire n3824_o;
  wire n3827_o;
  wire n3829_o;
  wire [2:0] n3830_o;
  wire n3832_o;
  wire [2:0] n3833_o;
  wire n3835_o;
  wire [1:0] n3836_o;
  wire n3838_o;
  wire n3839_o;
  wire n3840_o;
  wire [1:0] n3843_o;
  wire n3845_o;
  wire n3848_o;
  wire n3850_o;
  wire n3851_o;
  wire n3854_o;
  wire n3857_o;
  wire n3860_o;
  wire n3863_o;
  wire n3866_o;
  wire n3868_o;
  wire n3869_o;
  wire n3870_o;
  wire n3872_o;
  wire n3874_o;
  wire n3875_o;
  wire n3877_o;
  wire n3878_o;
  wire n3879_o;
  wire n3880_o;
  wire n3881_o;
  wire n3883_o;
  wire n3884_o;
  wire n3885_o;
  wire n3886_o;
  wire n3887_o;
  wire n3889_o;
  wire n3891_o;
  wire n3893_o;
  wire [1:0] n3894_o;
  wire n3896_o;
  wire [2:0] n3897_o;
  wire n3899_o;
  wire [3:0] n3900_o;
  wire n3902_o;
  wire [1:0] n3903_o;
  wire n3905_o;
  wire n3906_o;
  wire n3907_o;
  wire [1:0] n3908_o;
  wire n3910_o;
  wire n3911_o;
  wire n3913_o;
  wire n3914_o;
  wire n3915_o;
  wire n3916_o;
  wire n3917_o;
  wire [1:0] n3920_o;
  wire [1:0] n3921_o;
  wire [1:0] n3922_o;
  wire n3923_o;
  wire [1:0] n3924_o;
  wire n3926_o;
  wire n3927_o;
  wire n3928_o;
  wire n3930_o;
  wire n3931_o;
  wire n3932_o;
  wire n3933_o;
  wire n3934_o;
  wire [1:0] n3936_o;
  wire [1:0] n3938_o;
  wire n3939_o;
  wire n3942_o;
  wire n3945_o;
  wire n3948_o;
  wire n3951_o;
  wire n3953_o;
  wire n3954_o;
  wire n3955_o;
  wire n3957_o;
  wire n3960_o;
  wire n3962_o;
  wire n3964_o;
  wire n3966_o;
  wire n3968_o;
  wire [2:0] n3969_o;
  wire n3971_o;
  wire [2:0] n3972_o;
  wire n3974_o;
  wire [1:0] n3975_o;
  wire n3977_o;
  wire n3978_o;
  wire n3979_o;
  wire [2:0] n3982_o;
  wire n3984_o;
  wire n3987_o;
  wire n3989_o;
  wire n3990_o;
  wire n3993_o;
  wire n3996_o;
  wire n3999_o;
  wire n4002_o;
  wire n4004_o;
  wire n4006_o;
  wire n4008_o;
  wire n4010_o;
  wire n4011_o;
  wire n4012_o;
  wire n4014_o;
  wire n4016_o;
  wire n4017_o;
  wire n4019_o;
  wire n4020_o;
  wire n4021_o;
  wire n4023_o;
  wire n4024_o;
  wire n4025_o;
  wire n4027_o;
  wire n4029_o;
  wire n4031_o;
  wire n4033_o;
  wire n4034_o;
  wire [2:0] n4035_o;
  wire n4037_o;
  wire n4038_o;
  wire n4039_o;
  wire n4040_o;
  wire n4044_o;
  wire n4045_o;
  wire [1:0] n4048_o;
  wire n4050_o;
  wire n4051_o;
  wire n4052_o;
  wire [1:0] n4053_o;
  wire n4055_o;
  wire n4056_o;
  wire [2:0] n4057_o;
  wire n4059_o;
  wire [1:0] n4060_o;
  wire n4062_o;
  wire n4063_o;
  wire n4064_o;
  wire n4065_o;
  wire n4066_o;
  wire n4067_o;
  wire [1:0] n4068_o;
  wire n4070_o;
  wire [2:0] n4071_o;
  wire n4073_o;
  wire n4074_o;
  wire [3:0] n4075_o;
  wire n4077_o;
  wire n4078_o;
  wire n4079_o;
  wire n4080_o;
  wire n4082_o;
  wire n4083_o;
  wire [1:0] n4085_o;
  wire [2:0] n4086_o;
  wire n4088_o;
  wire [2:0] n4089_o;
  wire n4091_o;
  wire n4092_o;
  wire n4094_o;
  wire n4095_o;
  wire n4099_o;
  wire n4101_o;
  wire [2:0] n4102_o;
  wire n4104_o;
  wire n4108_o;
  wire n4109_o;
  wire n4110_o;
  wire n4112_o;
  wire n4113_o;
  wire n4114_o;
  wire n4117_o;
  wire n4118_o;
  wire n4119_o;
  wire n4120_o;
  wire [2:0] n4122_o;
  wire n4124_o;
  wire [2:0] n4125_o;
  wire n4127_o;
  wire n4128_o;
  wire [2:0] n4129_o;
  wire n4131_o;
  wire n4132_o;
  wire n4134_o;
  wire n4135_o;
  wire [6:0] n4138_o;
  wire n4139_o;
  wire n4140_o;
  wire n4141_o;
  wire n4142_o;
  wire [6:0] n4143_o;
  wire n4144_o;
  wire n4146_o;
  wire n4147_o;
  wire [1:0] n4151_o;
  wire n4152_o;
  wire n4153_o;
  wire [1:0] n4156_o;
  wire n4158_o;
  wire n4159_o;
  wire n4160_o;
  wire n4161_o;
  wire n4162_o;
  wire [6:0] n4164_o;
  wire [1:0] n4165_o;
  wire n4167_o;
  wire n4169_o;
  wire n4171_o;
  wire n4172_o;
  wire n4173_o;
  wire n4174_o;
  wire n4177_o;
  wire n4179_o;
  wire n4182_o;
  wire n4185_o;
  wire [1:0] n4186_o;
  wire n4188_o;
  wire n4190_o;
  wire n4192_o;
  wire n4194_o;
  wire [1:0] n4195_o;
  wire n4197_o;
  wire n4199_o;
  wire n4201_o;
  wire n4203_o;
  wire n4205_o;
  wire [6:0] n4206_o;
  wire [1:0] n4207_o;
  wire [1:0] n4208_o;
  wire n4210_o;
  wire n4213_o;
  wire n4215_o;
  wire n4217_o;
  wire n4219_o;
  wire n4220_o;
  wire n4221_o;
  wire n4222_o;
  wire n4223_o;
  wire n4224_o;
  wire n4225_o;
  wire n4226_o;
  wire n4227_o;
  wire [1:0] n4228_o;
  wire n4229_o;
  wire n4230_o;
  wire n4231_o;
  wire n4232_o;
  wire n4233_o;
  wire n4234_o;
  wire n4236_o;
  wire n4238_o;
  wire n4240_o;
  wire n4241_o;
  wire n4243_o;
  wire [6:0] n4244_o;
  wire n4245_o;
  wire [1:0] n4246_o;
  wire n4248_o;
  wire [2:0] n4249_o;
  wire n4251_o;
  wire n4252_o;
  wire [3:0] n4253_o;
  wire n4255_o;
  wire [1:0] n4256_o;
  wire n4258_o;
  wire n4259_o;
  wire n4260_o;
  wire n4262_o;
  wire n4263_o;
  wire n4264_o;
  wire n4265_o;
  wire n4267_o;
  wire n4269_o;
  wire n4270_o;
  wire n4271_o;
  wire n4274_o;
  wire n4275_o;
  wire n4276_o;
  wire n4277_o;
  wire [6:0] n4279_o;
  wire n4281_o;
  wire n4282_o;
  wire [1:0] n4283_o;
  wire n4285_o;
  wire n4286_o;
  wire n4287_o;
  wire n4288_o;
  wire n4291_o;
  wire [1:0] n4293_o;
  wire [6:0] n4295_o;
  wire n4299_o;
  wire n4302_o;
  wire n4303_o;
  wire n4304_o;
  wire n4305_o;
  wire n4306_o;
  wire n4307_o;
  wire n4308_o;
  wire n4309_o;
  wire [1:0] n4310_o;
  wire n4312_o;
  wire [2:0] n4313_o;
  wire n4315_o;
  wire n4316_o;
  wire [3:0] n4317_o;
  wire n4319_o;
  wire [1:0] n4320_o;
  wire n4322_o;
  wire n4323_o;
  wire n4324_o;
  wire n4325_o;
  wire n4326_o;
  wire n4328_o;
  wire n4330_o;
  wire n4331_o;
  wire n4332_o;
  wire n4333_o;
  wire n4334_o;
  wire n4336_o;
  wire n4338_o;
  wire n4339_o;
  wire n4340_o;
  wire n4341_o;
  wire n4344_o;
  wire n4345_o;
  wire n4346_o;
  wire n4347_o;
  wire [6:0] n4349_o;
  wire n4351_o;
  wire n4352_o;
  wire [1:0] n4353_o;
  wire n4355_o;
  wire n4356_o;
  wire n4357_o;
  wire n4358_o;
  wire n4359_o;
  wire n4361_o;
  wire n4362_o;
  wire [6:0] n4365_o;
  wire [1:0] n4367_o;
  wire n4370_o;
  wire n4373_o;
  wire n4374_o;
  wire n4375_o;
  wire [6:0] n4376_o;
  wire [1:0] n4377_o;
  wire n4379_o;
  wire n4380_o;
  wire n4381_o;
  wire n4384_o;
  wire [1:0] n4386_o;
  wire n4387_o;
  wire n4390_o;
  wire n4392_o;
  wire n4394_o;
  wire n4396_o;
  wire n4399_o;
  wire n4402_o;
  wire n4404_o;
  wire n4406_o;
  wire n4408_o;
  wire [6:0] n4409_o;
  wire [1:0] n4411_o;
  wire [1:0] n4412_o;
  wire n4414_o;
  wire n4416_o;
  wire n4417_o;
  wire n4419_o;
  wire n4421_o;
  wire n4423_o;
  wire n4425_o;
  wire n4426_o;
  wire n4427_o;
  wire n4429_o;
  wire n4430_o;
  wire n4432_o;
  wire n4433_o;
  wire [6:0] n4434_o;
  wire n4435_o;
  wire [2:0] n4436_o;
  wire n4438_o;
  wire [2:0] n4441_o;
  wire n4443_o;
  wire n4444_o;
  wire [1:0] n4445_o;
  wire n4447_o;
  wire n4448_o;
  wire [2:0] n4449_o;
  wire n4451_o;
  wire n4452_o;
  wire [3:0] n4453_o;
  wire n4455_o;
  wire n4456_o;
  wire n4458_o;
  wire n4459_o;
  wire [1:0] n4462_o;
  wire n4464_o;
  wire n4465_o;
  wire n4466_o;
  wire n4467_o;
  wire n4468_o;
  wire [6:0] n4470_o;
  wire n4471_o;
  wire [1:0] n4473_o;
  wire [1:0] n4474_o;
  wire n4475_o;
  wire n4478_o;
  wire n4481_o;
  wire n4484_o;
  wire n4487_o;
  wire n4488_o;
  wire n4489_o;
  wire n4490_o;
  wire n4491_o;
  wire n4492_o;
  wire [1:0] n4493_o;
  wire n4494_o;
  wire n4496_o;
  wire n4498_o;
  wire n4500_o;
  wire n4502_o;
  wire n4503_o;
  wire n4504_o;
  wire n4505_o;
  wire n4506_o;
  wire [6:0] n4507_o;
  wire [1:0] n4508_o;
  wire n4509_o;
  wire n4511_o;
  wire n4513_o;
  wire n4515_o;
  wire n4517_o;
  wire n4518_o;
  wire n4519_o;
  wire n4520_o;
  wire n4521_o;
  wire n4523_o;
  wire n4525_o;
  wire [6:0] n4526_o;
  wire [2:0] n4527_o;
  wire n4529_o;
  wire n4539_o;
  wire n4542_o;
  wire n4545_o;
  wire n4546_o;
  wire n4547_o;
  wire n4548_o;
  wire n4549_o;
  wire n4550_o;
  wire n4551_o;
  wire n4552_o;
  wire n4553_o;
  wire n4554_o;
  wire n4555_o;
  wire n4556_o;
  wire [6:0] n4558_o;
  wire [2:0] n4559_o;
  wire n4561_o;
  wire [2:0] n4562_o;
  wire n4564_o;
  wire [1:0] n4565_o;
  wire n4567_o;
  wire n4568_o;
  wire n4569_o;
  wire [1:0] n4574_o;
  wire n4576_o;
  wire n4579_o;
  wire n4581_o;
  wire n4582_o;
  wire n4585_o;
  wire n4588_o;
  wire n4591_o;
  wire n4594_o;
  wire n4597_o;
  wire n4599_o;
  wire n4600_o;
  wire n4601_o;
  wire n4603_o;
  wire n4605_o;
  wire n4607_o;
  wire n4609_o;
  wire [1:0] n4611_o;
  wire n4613_o;
  wire n4614_o;
  wire n4616_o;
  wire n4617_o;
  wire n4619_o;
  wire n4621_o;
  wire n4623_o;
  wire n4625_o;
  wire n4627_o;
  wire n4628_o;
  wire n4629_o;
  wire n4630_o;
  wire n4631_o;
  wire n4632_o;
  wire n4633_o;
  wire n4634_o;
  wire n4635_o;
  wire n4637_o;
  wire n4638_o;
  wire n4639_o;
  wire n4640_o;
  wire n4641_o;
  wire n4643_o;
  wire n4645_o;
  wire n4646_o;
  wire n4647_o;
  wire [1:0] n4649_o;
  wire [1:0] n4650_o;
  wire n4652_o;
  wire n4653_o;
  wire n4655_o;
  wire n4657_o;
  wire n4659_o;
  wire n4660_o;
  wire n4661_o;
  wire n4662_o;
  wire [2:0] n4663_o;
  wire n4664_o;
  wire n4665_o;
  wire n4666_o;
  wire n4667_o;
  wire n4668_o;
  wire n4669_o;
  wire n4670_o;
  wire [2:0] n4671_o;
  wire [2:0] n4672_o;
  wire n4673_o;
  wire n4675_o;
  wire n4677_o;
  wire n4679_o;
  wire n4681_o;
  wire n4682_o;
  wire [6:0] n4683_o;
  wire [1:0] n4684_o;
  wire [1:0] n4685_o;
  wire n4687_o;
  wire n4688_o;
  wire n4690_o;
  wire n4692_o;
  wire n4693_o;
  wire n4695_o;
  wire n4697_o;
  wire n4699_o;
  wire n4700_o;
  wire n4701_o;
  wire n4703_o;
  wire n4705_o;
  wire n4706_o;
  wire n4707_o;
  wire n4709_o;
  wire n4710_o;
  wire n4711_o;
  wire n4712_o;
  wire n4713_o;
  wire n4714_o;
  wire n4715_o;
  wire n4716_o;
  wire n4717_o;
  wire n4718_o;
  wire n4719_o;
  wire n4720_o;
  wire n4721_o;
  wire [2:0] n4722_o;
  wire [2:0] n4723_o;
  wire n4725_o;
  wire n4726_o;
  wire n4727_o;
  wire n4728_o;
  wire n4730_o;
  wire n4732_o;
  wire n4734_o;
  wire n4736_o;
  wire n4738_o;
  wire [6:0] n4739_o;
  wire [1:0] n4740_o;
  wire [1:0] n4741_o;
  wire n4743_o;
  wire n4744_o;
  wire n4745_o;
  wire n4747_o;
  wire n4748_o;
  wire n4750_o;
  wire n4752_o;
  wire n4754_o;
  wire n4756_o;
  wire n4757_o;
  wire n4758_o;
  wire n4760_o;
  wire n4761_o;
  wire n4762_o;
  wire n4763_o;
  wire n4764_o;
  wire n4765_o;
  wire n4766_o;
  wire n4767_o;
  wire n4768_o;
  wire n4769_o;
  wire n4770_o;
  wire n4771_o;
  wire n4772_o;
  wire n4773_o;
  wire n4774_o;
  wire n4775_o;
  wire n4776_o;
  wire n4777_o;
  wire n4778_o;
  wire n4779_o;
  wire n4780_o;
  wire n4781_o;
  wire n4782_o;
  wire n4783_o;
  wire n4784_o;
  wire n4785_o;
  wire n4786_o;
  wire n4787_o;
  wire n4788_o;
  wire n4789_o;
  wire n4790_o;
  wire n4791_o;
  wire n4792_o;
  wire n4793_o;
  wire n4794_o;
  wire n4795_o;
  wire n4796_o;
  wire n4797_o;
  wire n4799_o;
  wire n4801_o;
  wire n4803_o;
  wire n4805_o;
  wire n4807_o;
  wire n4809_o;
  wire n4811_o;
  wire n4812_o;
  wire n4814_o;
  wire [6:0] n4815_o;
  wire n4817_o;
  wire n4819_o;
  wire n4820_o;
  wire [4:0] n4821_o;
  wire n4823_o;
  wire [1:0] n4824_o;
  wire n4826_o;
  wire n4827_o;
  wire [1:0] n4828_o;
  wire n4830_o;
  wire [2:0] n4831_o;
  wire n4833_o;
  wire [2:0] n4834_o;
  wire n4836_o;
  wire [1:0] n4837_o;
  wire n4839_o;
  wire n4840_o;
  wire n4841_o;
  wire n4842_o;
  wire [1:0] n4843_o;
  wire n4845_o;
  wire [2:0] n4846_o;
  wire n4848_o;
  wire n4849_o;
  wire [3:0] n4850_o;
  wire n4852_o;
  wire [1:0] n4853_o;
  wire n4855_o;
  wire n4856_o;
  wire n4857_o;
  wire n4858_o;
  wire n4859_o;
  wire n4862_o;
  wire n4864_o;
  wire n4867_o;
  wire [1:0] n4869_o;
  wire n4871_o;
  wire [1:0] n4872_o;
  wire n4874_o;
  wire n4877_o;
  wire [1:0] n4879_o;
  wire n4882_o;
  wire n4885_o;
  wire n4887_o;
  wire n4888_o;
  wire n4890_o;
  wire n4892_o;
  wire n4894_o;
  wire n4896_o;
  wire n4899_o;
  wire n4902_o;
  wire n4905_o;
  wire n4907_o;
  wire n4909_o;
  wire [1:0] n4910_o;
  wire n4912_o;
  wire n4914_o;
  wire n4916_o;
  wire n4918_o;
  wire n4920_o;
  wire n4922_o;
  wire n4924_o;
  wire n4926_o;
  wire n4928_o;
  wire n4930_o;
  wire n4931_o;
  wire n4932_o;
  wire [1:0] n4933_o;
  wire n4935_o;
  wire n4936_o;
  wire [2:0] n4937_o;
  wire n4939_o;
  wire n4940_o;
  wire [3:0] n4941_o;
  wire n4943_o;
  wire n4944_o;
  wire n4945_o;
  wire [6:0] n4947_o;
  wire n4949_o;
  wire n4950_o;
  wire n4951_o;
  wire n4952_o;
  wire n4953_o;
  wire [1:0] n4956_o;
  wire n4958_o;
  wire n4959_o;
  wire n4960_o;
  wire n4961_o;
  wire n4962_o;
  wire [6:0] n4964_o;
  wire n4966_o;
  wire n4967_o;
  wire n4968_o;
  wire n4969_o;
  wire n4971_o;
  wire n4973_o;
  wire n4976_o;
  wire n4978_o;
  wire n4979_o;
  wire n4980_o;
  wire n4981_o;
  wire n4983_o;
  wire n4985_o;
  wire [1:0] n4987_o;
  wire n4988_o;
  wire n4989_o;
  wire n4990_o;
  wire [1:0] n4992_o;
  wire [1:0] n4993_o;
  wire n4994_o;
  wire n4996_o;
  wire n4999_o;
  wire n5002_o;
  wire n5005_o;
  wire n5008_o;
  wire [1:0] n5009_o;
  wire n5010_o;
  wire n5011_o;
  wire n5012_o;
  wire n5013_o;
  wire [1:0] n5014_o;
  wire [6:0] n5015_o;
  wire [6:0] n5016_o;
  wire n5018_o;
  wire n5020_o;
  wire n5021_o;
  wire n5023_o;
  wire n5024_o;
  wire n5026_o;
  wire n5027_o;
  wire n5029_o;
  wire n5030_o;
  wire n5032_o;
  wire n5033_o;
  wire n5035_o;
  wire n5036_o;
  wire n5038_o;
  wire n5039_o;
  wire n5041_o;
  wire n5042_o;
  wire n5044_o;
  wire n5045_o;
  wire n5047_o;
  wire n5048_o;
  wire n5050_o;
  wire n5051_o;
  wire n5053_o;
  wire n5054_o;
  wire n5056_o;
  wire n5057_o;
  wire n5059_o;
  wire n5060_o;
  wire n5062_o;
  wire n5063_o;
  wire n5071_o;
  wire n5074_o;
  wire n5077_o;
  wire n5078_o;
  wire n5079_o;
  wire n5080_o;
  wire n5081_o;
  wire n5082_o;
  wire n5083_o;
  wire n5084_o;
  wire n5085_o;
  wire [6:0] n5087_o;
  wire n5089_o;
  wire n5091_o;
  wire n5092_o;
  wire n5094_o;
  wire n5095_o;
  wire n5097_o;
  wire n5098_o;
  wire n5100_o;
  wire n5101_o;
  wire n5103_o;
  wire n5104_o;
  wire n5106_o;
  wire n5107_o;
  wire n5109_o;
  wire n5110_o;
  wire [1:0] n5117_o;
  wire n5119_o;
  wire n5122_o;
  wire n5125_o;
  wire n5126_o;
  wire n5127_o;
  wire n5128_o;
  wire n5129_o;
  wire [6:0] n5131_o;
  wire n5133_o;
  wire n5135_o;
  wire n5136_o;
  wire n5138_o;
  wire n5139_o;
  wire n5141_o;
  wire n5142_o;
  wire n5144_o;
  wire n5145_o;
  wire n5147_o;
  wire n5148_o;
  wire n5150_o;
  wire n5151_o;
  wire n5153_o;
  wire n5154_o;
  wire [1:0] n5157_o;
  wire n5160_o;
  wire n5163_o;
  wire n5166_o;
  wire n5169_o;
  wire n5170_o;
  wire n5171_o;
  wire n5172_o;
  wire n5173_o;
  wire n5175_o;
  wire n5177_o;
  wire n5178_o;
  wire n5180_o;
  wire n5181_o;
  wire n5183_o;
  wire n5184_o;
  wire n5186_o;
  wire n5187_o;
  wire n5189_o;
  wire n5190_o;
  wire n5192_o;
  wire n5193_o;
  wire n5195_o;
  wire n5196_o;
  wire [1:0] n5200_o;
  wire n5203_o;
  wire n5206_o;
  wire n5207_o;
  wire n5208_o;
  wire n5209_o;
  wire n5210_o;
  wire n5212_o;
  wire n5214_o;
  wire n5216_o;
  wire n5217_o;
  wire n5219_o;
  wire n5220_o;
  wire n5222_o;
  wire n5223_o;
  wire n5225_o;
  wire n5226_o;
  wire n5228_o;
  wire n5229_o;
  wire n5231_o;
  wire n5232_o;
  wire n5234_o;
  wire n5235_o;
  wire n5236_o;
  wire [5:0] n5240_o;
  wire n5241_o;
  wire n5242_o;
  wire [5:0] n5243_o;
  wire n5246_o;
  wire n5249_o;
  wire n5250_o;
  wire n5251_o;
  wire n5252_o;
  wire n5253_o;
  wire n5255_o;
  wire n5257_o;
  wire n5258_o;
  wire n5260_o;
  wire n5263_o;
  wire n5265_o;
  wire n5266_o;
  wire n5267_o;
  wire n5270_o;
  wire n5273_o;
  wire n5275_o;
  wire n5277_o;
  wire n5278_o;
  wire n5279_o;
  wire n5281_o;
  wire n5284_o;
  wire n5285_o;
  wire n5286_o;
  wire n5287_o;
  wire [1:0] n5289_o;
  wire n5291_o;
  wire [1:0] n5292_o;
  wire n5293_o;
  wire n5294_o;
  wire n5295_o;
  wire n5296_o;
  wire [1:0] n5297_o;
  wire [1:0] n5298_o;
  wire [6:0] n5300_o;
  wire n5301_o;
  wire n5302_o;
  wire n5305_o;
  wire n5308_o;
  wire n5309_o;
  wire n5310_o;
  wire n5311_o;
  wire n5312_o;
  wire n5314_o;
  wire n5315_o;
  wire n5317_o;
  wire n5319_o;
  wire n5320_o;
  wire [1:0] n5325_o;
  wire n5327_o;
  wire n5329_o;
  wire [1:0] n5330_o;
  wire n5331_o;
  wire n5332_o;
  wire n5333_o;
  wire n5334_o;
  wire [1:0] n5335_o;
  wire [1:0] n5336_o;
  wire [6:0] n5338_o;
  wire n5340_o;
  wire [1:0] n5345_o;
  wire n5347_o;
  wire [1:0] n5348_o;
  wire n5349_o;
  wire n5350_o;
  wire n5351_o;
  wire n5352_o;
  wire [1:0] n5353_o;
  wire [1:0] n5354_o;
  wire [6:0] n5356_o;
  wire n5358_o;
  wire [1:0] n5360_o;
  wire n5361_o;
  wire n5363_o;
  wire n5364_o;
  wire n5367_o;
  wire n5370_o;
  wire n5372_o;
  wire n5374_o;
  wire n5375_o;
  wire [11:0] n5376_o;
  wire n5378_o;
  wire n5380_o;
  wire n5382_o;
  wire n5383_o;
  wire n5384_o;
  wire n5385_o;
  wire [1:0] n5386_o;
  wire [1:0] n5387_o;
  wire n5388_o;
  wire n5389_o;
  wire n5393_o;
  wire n5395_o;
  wire n5397_o;
  wire [6:0] n5399_o;
  wire [1:0] n5401_o;
  wire n5402_o;
  wire n5405_o;
  wire n5408_o;
  wire [1:0] n5409_o;
  wire [1:0] n5410_o;
  wire [1:0] n5412_o;
  wire [6:0] n5413_o;
  wire [1:0] n5414_o;
  wire n5415_o;
  wire n5418_o;
  wire n5420_o;
  wire n5422_o;
  wire [1:0] n5423_o;
  wire [1:0] n5425_o;
  wire [6:0] n5426_o;
  wire n5428_o;
  wire n5430_o;
  wire n5431_o;
  wire [12:0] n5432_o;
  reg n5433_o;
  reg [1:0] n5438_o;
  reg [1:0] n5439_o;
  reg n5440_o;
  reg n5441_o;
  reg n5442_o;
  reg n5444_o;
  reg n5446_o;
  reg [5:0] n5447_o;
  reg n5448_o;
  reg n5451_o;
  reg n5453_o;
  reg n5456_o;
  reg n5458_o;
  reg n5462_o;
  reg n5464_o;
  wire n5465_o;
  reg n5466_o;
  wire n5467_o;
  reg n5468_o;
  wire n5469_o;
  reg n5470_o;
  wire n5471_o;
  reg n5472_o;
  wire n5473_o;
  wire n5474_o;
  wire n5475_o;
  reg n5476_o;
  wire n5477_o;
  wire n5478_o;
  wire n5479_o;
  reg n5480_o;
  wire n5481_o;
  reg n5482_o;
  wire n5483_o;
  reg n5484_o;
  wire [1:0] n5485_o;
  reg [1:0] n5486_o;
  wire [1:0] n5487_o;
  reg [1:0] n5488_o;
  wire n5489_o;
  wire n5490_o;
  wire n5491_o;
  wire n5492_o;
  reg n5493_o;
  wire n5494_o;
  wire n5495_o;
  wire n5496_o;
  wire n5497_o;
  reg n5498_o;
  wire n5499_o;
  reg n5500_o;
  reg n5502_o;
  reg n5504_o;
  reg [1:0] n5506_o;
  reg n5508_o;
  reg [6:0] n5509_o;
  wire n5510_o;
  wire [1:0] n5511_o;
  wire [1:0] n5512_o;
  wire n5513_o;
  wire n5514_o;
  wire n5515_o;
  wire n5517_o;
  wire n5519_o;
  wire n5521_o;
  wire n5523_o;
  wire [5:0] n5524_o;
  wire n5525_o;
  wire n5526_o;
  wire n5528_o;
  wire n5530_o;
  wire n5532_o;
  wire n5533_o;
  wire n5535_o;
  wire n5537_o;
  wire [1:0] n5538_o;
  wire [3:0] n5539_o;
  wire [1:0] n5540_o;
  wire n5541_o;
  wire n5542_o;
  wire n5543_o;
  wire n5544_o;
  wire n5545_o;
  wire n5546_o;
  wire n5547_o;
  wire n5548_o;
  wire n5549_o;
  wire n5550_o;
  wire n5551_o;
  wire n5552_o;
  wire n5553_o;
  wire n5554_o;
  wire n5555_o;
  wire n5556_o;
  wire n5557_o;
  wire n5558_o;
  wire n5559_o;
  wire [3:0] n5560_o;
  wire [3:0] n5561_o;
  wire n5562_o;
  wire [1:0] n5563_o;
  wire n5564_o;
  wire n5565_o;
  wire [2:0] n5566_o;
  wire n5568_o;
  wire n5570_o;
  wire [2:0] n5572_o;
  wire [6:0] n5573_o;
  wire n5575_o;
  wire [6:0] n5576_o;
  reg n5577_o;
  reg [1:0] n5578_o;
  reg [1:0] n5579_o;
  reg n5580_o;
  reg n5581_o;
  reg n5583_o;
  reg n5584_o;
  reg n5586_o;
  reg n5588_o;
  reg n5590_o;
  reg n5592_o;
  reg n5594_o;
  reg n5596_o;
  reg n5598_o;
  reg n5600_o;
  reg [5:0] n5601_o;
  reg n5603_o;
  reg n5604_o;
  reg n5606_o;
  reg n5608_o;
  reg n5610_o;
  reg n5612_o;
  reg n5614_o;
  reg n5616_o;
  reg n5618_o;
  wire n5619_o;
  reg n5620_o;
  wire n5621_o;
  reg n5622_o;
  wire n5623_o;
  reg n5624_o;
  wire n5625_o;
  reg n5626_o;
  wire n5627_o;
  reg n5628_o;
  wire n5629_o;
  reg n5630_o;
  wire n5631_o;
  reg n5632_o;
  wire n5633_o;
  reg n5634_o;
  wire n5635_o;
  wire n5636_o;
  wire n5637_o;
  reg n5638_o;
  wire n5639_o;
  wire n5640_o;
  wire n5641_o;
  reg n5642_o;
  wire n5643_o;
  reg n5644_o;
  wire n5645_o;
  reg n5646_o;
  wire n5647_o;
  wire n5648_o;
  reg n5649_o;
  wire n5650_o;
  wire n5651_o;
  reg n5652_o;
  wire n5653_o;
  reg n5654_o;
  wire n5655_o;
  reg n5656_o;
  wire n5657_o;
  reg n5658_o;
  wire n5659_o;
  reg n5660_o;
  wire [3:0] n5661_o;
  reg [3:0] n5662_o;
  reg [1:0] n5663_o;
  reg [1:0] n5664_o;
  wire n5665_o;
  reg n5666_o;
  wire n5667_o;
  reg n5668_o;
  wire n5669_o;
  reg n5670_o;
  reg n5671_o;
  wire n5672_o;
  reg n5673_o;
  reg n5675_o;
  wire n5676_o;
  reg n5678_o;
  wire n5679_o;
  reg n5681_o;
  reg n5683_o;
  reg n5685_o;
  reg n5687_o;
  reg n5689_o;
  reg n5691_o;
  reg n5693_o;
  reg n5695_o;
  reg n5697_o;
  wire [1:0] n5698_o;
  reg [1:0] n5700_o;
  wire n5701_o;
  reg n5703_o;
  reg n5705_o;
  reg [6:0] n5706_o;
  wire n5707_o;
  wire [1:0] n5708_o;
  wire [1:0] n5709_o;
  wire n5710_o;
  wire n5711_o;
  wire n5713_o;
  wire n5714_o;
  wire n5716_o;
  wire n5718_o;
  wire n5719_o;
  wire n5720_o;
  wire n5721_o;
  wire n5723_o;
  wire n5725_o;
  wire n5727_o;
  wire n5728_o;
  wire [5:0] n5729_o;
  wire n5731_o;
  wire n5732_o;
  wire n5733_o;
  wire n5735_o;
  wire n5737_o;
  wire n5739_o;
  wire n5740_o;
  wire n5742_o;
  wire n5743_o;
  wire [3:0] n5744_o;
  wire [9:0] n5745_o;
  wire [4:0] n5746_o;
  wire [1:0] n5747_o;
  wire n5748_o;
  wire n5749_o;
  wire n5750_o;
  wire n5751_o;
  wire n5752_o;
  wire n5753_o;
  wire n5754_o;
  wire n5755_o;
  wire n5756_o;
  wire n5757_o;
  wire n5758_o;
  wire n5759_o;
  wire n5760_o;
  wire n5761_o;
  wire n5762_o;
  wire n5763_o;
  wire n5764_o;
  wire n5765_o;
  wire [2:0] n5766_o;
  wire n5767_o;
  wire [2:0] n5768_o;
  wire [2:0] n5769_o;
  wire n5770_o;
  wire n5771_o;
  wire [4:0] n5772_o;
  wire [4:0] n5773_o;
  wire [4:0] n5774_o;
  wire n5775_o;
  wire n5776_o;
  wire [3:0] n5777_o;
  wire [3:0] n5778_o;
  wire [3:0] n5779_o;
  wire n5780_o;
  wire [4:0] n5781_o;
  wire [4:0] n5782_o;
  wire n5783_o;
  wire n5784_o;
  wire n5785_o;
  wire n5786_o;
  wire n5787_o;
  wire [1:0] n5788_o;
  wire [1:0] n5789_o;
  wire [1:0] n5790_o;
  wire [1:0] n5791_o;
  wire [2:0] n5792_o;
  wire n5793_o;
  wire [1:0] n5795_o;
  wire [1:0] n5797_o;
  wire n5798_o;
  wire n5800_o;
  wire n5802_o;
  wire n5804_o;
  wire n5806_o;
  wire n5808_o;
  wire n5810_o;
  wire [1:0] n5811_o;
  wire [1:0] n5813_o;
  wire n5814_o;
  wire n5815_o;
  wire n5816_o;
  wire [6:0] n5817_o;
  wire n5819_o;
  wire [1:0] n5820_o;
  wire n5822_o;
  wire [2:0] n5823_o;
  wire n5825_o;
  wire n5829_o;
  wire n5830_o;
  wire n5831_o;
  wire [6:0] n5833_o;
  wire [2:0] n5834_o;
  wire n5836_o;
  wire [1:0] n5837_o;
  wire n5839_o;
  wire [2:0] n5840_o;
  wire n5842_o;
  wire n5843_o;
  wire n5844_o;
  wire n5845_o;
  wire [1:0] n5846_o;
  wire n5848_o;
  wire n5849_o;
  wire n5851_o;
  wire n5852_o;
  wire [6:0] n5854_o;
  wire [1:0] n5856_o;
  wire [1:0] n5857_o;
  wire n5858_o;
  wire n5859_o;
  wire n5860_o;
  wire n5861_o;
  wire n5864_o;
  wire n5867_o;
  wire [1:0] n5868_o;
  wire n5871_o;
  wire n5873_o;
  wire n5875_o;
  wire n5876_o;
  wire n5877_o;
  wire [2:0] n5878_o;
  wire n5880_o;
  wire [1:0] n5881_o;
  wire n5883_o;
  wire n5884_o;
  wire n5886_o;
  wire n5888_o;
  wire n5889_o;
  wire n5890_o;
  wire n5891_o;
  wire n5893_o;
  wire [1:0] n5894_o;
  wire n5896_o;
  wire n5899_o;
  wire n5900_o;
  wire [1:0] n5902_o;
  wire n5905_o;
  wire n5908_o;
  wire n5911_o;
  wire n5914_o;
  wire n5916_o;
  wire n5918_o;
  wire n5919_o;
  wire [1:0] n5920_o;
  wire n5921_o;
  wire n5923_o;
  wire n5924_o;
  wire n5926_o;
  wire n5927_o;
  wire n5929_o;
  wire n5930_o;
  wire n5932_o;
  wire n5934_o;
  wire n5935_o;
  wire n5936_o;
  wire [1:0] n5937_o;
  wire [1:0] n5938_o;
  wire n5940_o;
  wire n5942_o;
  wire n5944_o;
  wire n5946_o;
  wire n5948_o;
  wire n5950_o;
  wire n5952_o;
  wire n5953_o;
  wire n5955_o;
  wire n5957_o;
  wire [6:0] n5958_o;
  wire [4:0] n5959_o;
  wire n5961_o;
  wire [2:0] n5962_o;
  wire n5964_o;
  wire [1:0] n5965_o;
  wire n5967_o;
  wire n5968_o;
  wire n5969_o;
  wire [2:0] n5970_o;
  wire n5972_o;
  wire n5974_o;
  wire n5975_o;
  wire n5976_o;
  wire n5978_o;
  wire n5979_o;
  wire [1:0] n5983_o;
  wire n5985_o;
  wire n5988_o;
  wire n5991_o;
  wire n5994_o;
  wire n5997_o;
  wire n6000_o;
  wire n6002_o;
  wire n6004_o;
  wire [1:0] n6005_o;
  wire [1:0] n6007_o;
  wire n6009_o;
  wire n6011_o;
  wire n6012_o;
  wire [1:0] n6013_o;
  wire [1:0] n6014_o;
  wire n6016_o;
  wire n6017_o;
  wire n6018_o;
  wire n6020_o;
  wire n6021_o;
  wire n6022_o;
  wire n6023_o;
  wire n6024_o;
  wire n6026_o;
  wire n6027_o;
  wire n6028_o;
  wire n6029_o;
  wire [1:0] n6031_o;
  wire n6033_o;
  wire n6035_o;
  wire n6036_o;
  wire [6:0] n6037_o;
  wire n6039_o;
  wire n6041_o;
  wire [3:0] n6042_o;
  wire n6044_o;
  wire [7:0] n6046_o;
  wire n6048_o;
  wire [7:0] n6050_o;
  wire n6052_o;
  wire [1:0] n6054_o;
  wire n6057_o;
  wire [6:0] n6060_o;
  wire [1:0] n6061_o;
  wire n6063_o;
  wire n6064_o;
  wire [6:0] n6066_o;
  wire [7:0] n6067_o;
  wire n6069_o;
  wire [7:0] n6071_o;
  wire n6073_o;
  wire [1:0] n6075_o;
  wire [1:0] n6076_o;
  wire n6077_o;
  wire [1:0] n6078_o;
  wire n6080_o;
  wire n6082_o;
  wire n6083_o;
  wire n6084_o;
  wire n6085_o;
  wire n6086_o;
  wire n6087_o;
  wire [6:0] n6089_o;
  wire [1:0] n6090_o;
  wire n6091_o;
  wire n6093_o;
  wire n6094_o;
  wire n6095_o;
  wire n6096_o;
  wire n6097_o;
  wire n6098_o;
  wire [6:0] n6099_o;
  wire n6101_o;
  wire n6102_o;
  wire n6103_o;
  wire [1:0] n6108_o;
  wire n6111_o;
  wire n6114_o;
  wire n6117_o;
  wire [1:0] n6118_o;
  wire [1:0] n6120_o;
  wire n6122_o;
  wire n6124_o;
  wire [1:0] n6125_o;
  wire n6127_o;
  wire [2:0] n6128_o;
  wire n6130_o;
  wire n6132_o;
  wire [3:0] n6133_o;
  wire n6135_o;
  wire [1:0] n6136_o;
  wire n6138_o;
  wire n6139_o;
  wire n6140_o;
  wire [1:0] n6141_o;
  wire n6143_o;
  wire n6146_o;
  wire n6148_o;
  wire n6149_o;
  wire [1:0] n6150_o;
  wire n6152_o;
  wire n6153_o;
  wire n6154_o;
  wire [1:0] n6156_o;
  wire [6:0] n6158_o;
  wire n6159_o;
  wire n6160_o;
  wire n6161_o;
  wire n6164_o;
  wire [1:0] n6165_o;
  wire n6167_o;
  wire n6168_o;
  wire n6169_o;
  wire n6172_o;
  wire [1:0] n6174_o;
  wire n6175_o;
  wire n6177_o;
  wire n6180_o;
  wire n6182_o;
  wire n6185_o;
  wire n6188_o;
  wire n6191_o;
  wire n6193_o;
  wire n6194_o;
  wire n6195_o;
  wire [1:0] n6196_o;
  wire n6198_o;
  wire n6199_o;
  wire [1:0] n6200_o;
  wire n6202_o;
  wire [1:0] n6206_o;
  wire n6208_o;
  wire [1:0] n6209_o;
  wire n6211_o;
  wire n6212_o;
  wire [1:0] n6215_o;
  wire n6217_o;
  wire [1:0] n6222_o;
  wire n6224_o;
  wire n6226_o;
  wire n6227_o;
  wire n6228_o;
  wire [1:0] n6229_o;
  wire n6231_o;
  wire [1:0] n6234_o;
  wire n6238_o;
  wire n6239_o;
  wire n6240_o;
  wire n6241_o;
  wire [6:0] n6243_o;
  wire n6245_o;
  wire [6:0] n6247_o;
  wire [1:0] n6248_o;
  wire n6251_o;
  wire n6254_o;
  wire n6255_o;
  wire n6257_o;
  wire n6259_o;
  wire n6261_o;
  wire [6:0] n6262_o;
  wire [1:0] n6263_o;
  wire n6264_o;
  wire n6266_o;
  wire n6269_o;
  wire n6271_o;
  wire n6272_o;
  wire n6275_o;
  wire n6278_o;
  wire n6280_o;
  wire n6281_o;
  wire n6282_o;
  wire n6284_o;
  wire [1:0] n6285_o;
  wire n6287_o;
  wire n6289_o;
  wire [1:0] n6291_o;
  wire [6:0] n6292_o;
  wire [1:0] n6293_o;
  wire [1:0] n6294_o;
  wire n6296_o;
  wire n6298_o;
  wire n6300_o;
  wire n6301_o;
  wire n6303_o;
  wire n6305_o;
  wire n6308_o;
  wire n6309_o;
  wire n6310_o;
  wire n6311_o;
  wire n6312_o;
  wire n6313_o;
  wire n6314_o;
  wire n6315_o;
  wire n6316_o;
  wire n6318_o;
  wire n6320_o;
  wire n6322_o;
  wire n6324_o;
  wire [1:0] n6326_o;
  wire [6:0] n6327_o;
  wire [1:0] n6328_o;
  wire n6330_o;
  wire n6331_o;
  wire n6332_o;
  wire [2:0] n6333_o;
  wire n6335_o;
  wire n6336_o;
  wire [3:0] n6337_o;
  wire n6339_o;
  wire [1:0] n6340_o;
  wire n6342_o;
  wire n6343_o;
  wire n6344_o;
  wire n6345_o;
  wire [1:0] n6346_o;
  wire n6348_o;
  wire n6349_o;
  wire [2:0] n6350_o;
  wire n6352_o;
  wire [1:0] n6353_o;
  wire n6355_o;
  wire n6356_o;
  wire n6357_o;
  wire n6358_o;
  wire n6359_o;
  wire n6363_o;
  wire n6366_o;
  wire n6369_o;
  wire n6371_o;
  wire [1:0] n6372_o;
  wire [1:0] n6373_o;
  wire n6375_o;
  wire n6377_o;
  wire n6379_o;
  wire n6380_o;
  wire n6381_o;
  wire n6382_o;
  wire n6384_o;
  wire n6386_o;
  wire n6387_o;
  wire n6388_o;
  wire n6389_o;
  wire n6390_o;
  wire n6392_o;
  wire n6393_o;
  wire n6394_o;
  wire n6396_o;
  wire n6398_o;
  wire n6400_o;
  wire n6402_o;
  wire n6404_o;
  wire [1:0] n6406_o;
  wire [6:0] n6407_o;
  wire [1:0] n6408_o;
  wire [1:0] n6409_o;
  wire n6410_o;
  wire n6412_o;
  wire n6414_o;
  wire n6415_o;
  wire n6416_o;
  wire n6417_o;
  wire n6418_o;
  wire n6419_o;
  wire n6421_o;
  wire n6423_o;
  wire n6425_o;
  wire n6426_o;
  wire n6427_o;
  wire n6428_o;
  wire n6429_o;
  wire n6430_o;
  wire n6431_o;
  wire n6432_o;
  wire n6433_o;
  wire n6435_o;
  wire n6437_o;
  wire n6439_o;
  wire n6441_o;
  wire n6442_o;
  wire [1:0] n6444_o;
  wire [6:0] n6445_o;
  wire n6447_o;
  wire [5:0] n6448_o;
  wire n6450_o;
  wire n6451_o;
  wire n6452_o;
  wire [1:0] n6453_o;
  wire n6455_o;
  wire n6456_o;
  wire [3:0] n6457_o;
  wire n6459_o;
  wire [1:0] n6460_o;
  wire n6462_o;
  wire n6463_o;
  wire n6464_o;
  wire n6465_o;
  wire [2:0] n6466_o;
  wire n6468_o;
  wire [1:0] n6469_o;
  wire n6471_o;
  wire n6472_o;
  wire n6473_o;
  wire n6474_o;
  wire n6475_o;
  wire n6477_o;
  wire n6478_o;
  wire n6480_o;
  wire n6481_o;
  wire [1:0] n6482_o;
  wire n6484_o;
  wire n6485_o;
  wire n6486_o;
  wire [1:0] n6488_o;
  wire n6490_o;
  wire n6493_o;
  wire n6497_o;
  wire n6500_o;
  wire n6501_o;
  wire [1:0] n6502_o;
  wire n6504_o;
  wire n6505_o;
  wire n6508_o;
  wire n6511_o;
  wire n6512_o;
  wire n6514_o;
  wire n6517_o;
  wire n6519_o;
  wire n6521_o;
  wire n6523_o;
  wire n6525_o;
  wire n6526_o;
  wire n6527_o;
  wire n6529_o;
  wire n6530_o;
  wire n6532_o;
  wire n6534_o;
  wire n6536_o;
  wire n6538_o;
  wire n6541_o;
  wire n6544_o;
  wire n6547_o;
  wire n6549_o;
  wire n6551_o;
  wire n6553_o;
  wire n6555_o;
  wire n6557_o;
  wire n6559_o;
  wire n6561_o;
  wire n6563_o;
  wire n6564_o;
  wire n6566_o;
  wire [1:0] n6567_o;
  wire n6569_o;
  wire [3:0] n6570_o;
  wire n6572_o;
  wire [1:0] n6573_o;
  wire n6575_o;
  wire n6576_o;
  wire n6577_o;
  wire n6578_o;
  wire [1:0] n6581_o;
  wire n6583_o;
  wire n6585_o;
  wire n6588_o;
  wire n6590_o;
  wire n6593_o;
  wire n6596_o;
  wire n6599_o;
  wire n6601_o;
  wire n6603_o;
  wire n6605_o;
  wire n6607_o;
  wire n6609_o;
  wire n6612_o;
  wire n6615_o;
  wire n6618_o;
  wire n6619_o;
  wire n6620_o;
  wire n6622_o;
  wire n6624_o;
  wire n6625_o;
  wire [2:0] n6626_o;
  wire n6628_o;
  wire [2:0] n6630_o;
  wire n6632_o;
  wire n6634_o;
  wire [1:0] n6638_o;
  wire n6639_o;
  wire n6640_o;
  wire n6641_o;
  wire n6642_o;
  wire n6643_o;
  wire n6644_o;
  wire [6:0] n6646_o;
  wire [2:0] n6649_o;
  wire n6651_o;
  wire [1:0] n6652_o;
  wire n6654_o;
  wire n6655_o;
  wire n6659_o;
  wire n6662_o;
  wire n6665_o;
  wire n6668_o;
  wire n6670_o;
  wire n6671_o;
  wire n6673_o;
  wire n6675_o;
  wire n6677_o;
  wire n6679_o;
  wire n6680_o;
  wire n6681_o;
  wire n6682_o;
  wire n6683_o;
  wire n6684_o;
  wire n6685_o;
  wire n6686_o;
  wire n6687_o;
  wire n6689_o;
  wire n6691_o;
  wire n6693_o;
  wire n6694_o;
  wire [5:0] n6695_o;
  wire n6697_o;
  wire [3:0] n6698_o;
  wire n6700_o;
  wire [1:0] n6701_o;
  wire n6703_o;
  wire n6704_o;
  wire n6705_o;
  wire n6710_o;
  wire n6713_o;
  wire n6716_o;
  wire n6719_o;
  wire n6720_o;
  wire n6721_o;
  wire n6723_o;
  wire n6724_o;
  wire n6725_o;
  wire n6726_o;
  wire n6727_o;
  wire n6728_o;
  wire n6729_o;
  wire n6730_o;
  wire n6731_o;
  wire n6732_o;
  wire n6733_o;
  wire n6734_o;
  wire n6735_o;
  wire [1:0] n6736_o;
  wire n6737_o;
  wire n6739_o;
  wire n6740_o;
  wire n6741_o;
  wire n6743_o;
  wire n6744_o;
  wire n6745_o;
  wire [1:0] n6746_o;
  wire n6748_o;
  wire n6750_o;
  wire n6752_o;
  wire n6754_o;
  wire n6755_o;
  wire n6756_o;
  wire n6757_o;
  wire n6759_o;
  wire n6760_o;
  wire n6761_o;
  wire n6762_o;
  wire n6763_o;
  wire n6764_o;
  wire n6765_o;
  wire n6766_o;
  wire [1:0] n6767_o;
  wire n6768_o;
  wire n6770_o;
  wire n6771_o;
  wire n6772_o;
  wire n6774_o;
  wire n6776_o;
  wire [6:0] n6777_o;
  wire n6779_o;
  wire [1:0] n6780_o;
  wire n6782_o;
  wire [2:0] n6783_o;
  wire n6785_o;
  wire n6787_o;
  wire [3:0] n6788_o;
  wire n6790_o;
  wire [1:0] n6791_o;
  wire n6793_o;
  wire n6794_o;
  wire n6795_o;
  wire [1:0] n6796_o;
  wire n6798_o;
  wire n6801_o;
  wire n6803_o;
  wire n6804_o;
  wire [1:0] n6805_o;
  wire n6807_o;
  wire n6808_o;
  wire n6809_o;
  wire n6813_o;
  wire n6815_o;
  wire [1:0] n6817_o;
  wire n6819_o;
  wire n6820_o;
  wire n6821_o;
  wire n6824_o;
  wire [1:0] n6827_o;
  wire [1:0] n6829_o;
  wire n6831_o;
  wire n6834_o;
  wire n6836_o;
  wire n6839_o;
  wire n6842_o;
  wire n6845_o;
  wire n6847_o;
  wire n6849_o;
  wire n6851_o;
  wire n6852_o;
  wire [1:0] n6853_o;
  wire n6855_o;
  wire n6856_o;
  wire [1:0] n6857_o;
  wire n6859_o;
  wire [3:0] n6862_o;
  wire n6864_o;
  wire [4:0] n6865_o;
  wire n6867_o;
  wire n6868_o;
  wire n6872_o;
  wire n6873_o;
  wire n6874_o;
  wire n6877_o;
  wire n6880_o;
  wire [1:0] n6882_o;
  wire n6885_o;
  wire [1:0] n6887_o;
  wire n6888_o;
  wire n6890_o;
  wire n6892_o;
  wire n6894_o;
  wire n6897_o;
  wire n6900_o;
  wire n6901_o;
  wire n6902_o;
  wire n6903_o;
  wire n6904_o;
  wire n6905_o;
  wire n6906_o;
  wire [1:0] n6907_o;
  wire [1:0] n6908_o;
  wire n6910_o;
  wire n6912_o;
  wire n6914_o;
  wire n6916_o;
  wire n6918_o;
  wire n6921_o;
  wire n6922_o;
  wire n6923_o;
  wire n6924_o;
  wire n6925_o;
  wire n6926_o;
  wire n6927_o;
  wire n6929_o;
  wire n6931_o;
  wire [1:0] n6932_o;
  wire n6934_o;
  wire n6935_o;
  wire n6936_o;
  wire [2:0] n6937_o;
  wire n6939_o;
  wire n6940_o;
  wire [3:0] n6941_o;
  wire n6943_o;
  wire [1:0] n6944_o;
  wire n6946_o;
  wire n6947_o;
  wire n6948_o;
  wire n6949_o;
  wire [1:0] n6950_o;
  wire n6952_o;
  wire n6953_o;
  wire [2:0] n6954_o;
  wire n6956_o;
  wire [1:0] n6957_o;
  wire n6959_o;
  wire n6960_o;
  wire n6961_o;
  wire n6962_o;
  wire n6963_o;
  wire n6967_o;
  wire n6970_o;
  wire n6973_o;
  wire n6975_o;
  wire [1:0] n6976_o;
  wire [1:0] n6977_o;
  wire n6979_o;
  wire n6981_o;
  wire n6983_o;
  wire n6984_o;
  wire n6985_o;
  wire n6987_o;
  wire n6989_o;
  wire n6990_o;
  wire n6991_o;
  wire n6992_o;
  wire n6993_o;
  wire n6994_o;
  wire n6995_o;
  wire n6997_o;
  wire n6999_o;
  wire n7001_o;
  wire [1:0] n7002_o;
  wire [1:0] n7003_o;
  wire n7005_o;
  wire n7007_o;
  wire n7009_o;
  wire n7011_o;
  wire n7012_o;
  wire n7013_o;
  wire n7014_o;
  wire n7016_o;
  wire n7018_o;
  wire n7020_o;
  wire n7021_o;
  wire n7022_o;
  wire n7023_o;
  wire n7024_o;
  wire n7025_o;
  wire n7026_o;
  wire n7028_o;
  wire n7030_o;
  wire n7032_o;
  wire n7034_o;
  wire n7036_o;
  wire n7038_o;
  wire n7040_o;
  wire [1:0] n7041_o;
  wire n7043_o;
  wire n7044_o;
  wire n7045_o;
  wire [1:0] n7046_o;
  wire n7048_o;
  wire [2:0] n7049_o;
  wire n7051_o;
  wire [1:0] n7052_o;
  wire n7054_o;
  wire n7055_o;
  wire n7056_o;
  wire [1:0] n7058_o;
  wire [1:0] n7061_o;
  wire n7064_o;
  wire [1:0] n7065_o;
  wire n7068_o;
  wire n7071_o;
  wire n7074_o;
  wire n7076_o;
  wire n7078_o;
  wire n7079_o;
  wire n7080_o;
  wire n7082_o;
  wire n7084_o;
  wire [1:0] n7085_o;
  wire n7087_o;
  wire [2:0] n7088_o;
  wire n7090_o;
  wire n7091_o;
  wire [2:0] n7092_o;
  wire n7094_o;
  wire n7095_o;
  wire [2:0] n7096_o;
  wire n7098_o;
  wire [2:0] n7099_o;
  wire n7101_o;
  wire n7102_o;
  wire [2:0] n7103_o;
  wire n7105_o;
  wire n7106_o;
  wire [2:0] n7107_o;
  wire n7109_o;
  wire [1:0] n7110_o;
  wire n7112_o;
  wire n7113_o;
  wire n7114_o;
  wire n7115_o;
  wire n7116_o;
  wire [1:0] n7117_o;
  wire n7119_o;
  wire [2:0] n7120_o;
  wire n7122_o;
  wire n7123_o;
  wire [2:0] n7124_o;
  wire n7126_o;
  wire n7127_o;
  wire [2:0] n7128_o;
  wire n7130_o;
  wire [2:0] n7131_o;
  wire n7133_o;
  wire n7134_o;
  wire [2:0] n7135_o;
  wire n7137_o;
  wire n7138_o;
  wire [3:0] n7139_o;
  wire n7141_o;
  wire n7142_o;
  wire n7143_o;
  wire n7144_o;
  wire n7147_o;
  wire n7148_o;
  wire n7149_o;
  wire n7150_o;
  wire [6:0] n7152_o;
  wire n7154_o;
  wire n7155_o;
  wire n7156_o;
  wire n7157_o;
  wire n7160_o;
  wire [2:0] n7161_o;
  wire n7163_o;
  wire n7166_o;
  wire [2:0] n7167_o;
  wire n7169_o;
  wire [2:0] n7170_o;
  wire n7172_o;
  wire n7173_o;
  wire [2:0] n7174_o;
  wire n7176_o;
  wire n7177_o;
  wire [2:0] n7178_o;
  wire n7180_o;
  wire n7181_o;
  wire n7184_o;
  wire [2:0] n7185_o;
  wire n7187_o;
  wire [2:0] n7188_o;
  wire n7190_o;
  wire n7191_o;
  wire [2:0] n7192_o;
  wire n7194_o;
  wire n7195_o;
  wire n7198_o;
  wire [1:0] n7199_o;
  wire n7201_o;
  wire [2:0] n7202_o;
  wire n7204_o;
  wire n7206_o;
  wire n7207_o;
  wire [1:0] n7210_o;
  wire n7213_o;
  wire n7216_o;
  wire n7217_o;
  wire n7218_o;
  wire n7219_o;
  wire n7221_o;
  wire n7223_o;
  wire n7225_o;
  wire n7226_o;
  wire n7227_o;
  wire [1:0] n7229_o;
  wire n7230_o;
  wire [1:0] n7234_o;
  wire n7236_o;
  wire n7238_o;
  wire n7239_o;
  wire n7240_o;
  wire n7241_o;
  wire [6:0] n7243_o;
  wire [2:0] n7244_o;
  wire n7246_o;
  wire n7249_o;
  wire n7252_o;
  wire [2:0] n7253_o;
  wire n7255_o;
  wire [2:0] n7256_o;
  wire n7258_o;
  wire n7259_o;
  wire [2:0] n7260_o;
  wire n7262_o;
  wire n7263_o;
  wire n7265_o;
  wire n7267_o;
  wire n7269_o;
  wire n7270_o;
  wire [1:0] n7271_o;
  wire n7273_o;
  wire n7276_o;
  wire n7278_o;
  wire n7280_o;
  wire n7282_o;
  wire n7284_o;
  wire n7287_o;
  wire n7290_o;
  wire n7291_o;
  wire n7292_o;
  wire n7293_o;
  wire n7294_o;
  wire n7295_o;
  wire n7296_o;
  wire n7297_o;
  wire n7298_o;
  wire [1:0] n7299_o;
  wire n7301_o;
  wire n7303_o;
  wire [1:0] n7305_o;
  wire [6:0] n7306_o;
  wire n7307_o;
  wire [1:0] n7308_o;
  wire n7309_o;
  wire n7311_o;
  wire n7313_o;
  wire n7315_o;
  wire n7317_o;
  wire n7319_o;
  wire n7320_o;
  wire n7321_o;
  wire n7322_o;
  wire n7324_o;
  wire n7325_o;
  wire n7326_o;
  wire n7327_o;
  wire n7328_o;
  wire n7329_o;
  wire n7330_o;
  wire n7331_o;
  wire n7332_o;
  wire n7333_o;
  wire n7335_o;
  wire [1:0] n7337_o;
  wire n7339_o;
  wire [6:0] n7340_o;
  wire n7346_o;
  wire [1:0] n7347_o;
  wire n7350_o;
  wire n7352_o;
  wire n7354_o;
  wire n7356_o;
  wire n7358_o;
  wire n7360_o;
  wire n7362_o;
  wire n7363_o;
  wire n7365_o;
  wire n7367_o;
  wire n7369_o;
  wire n7370_o;
  wire n7371_o;
  wire n7372_o;
  wire n7373_o;
  wire n7374_o;
  wire n7375_o;
  wire n7376_o;
  wire n7377_o;
  wire n7379_o;
  wire n7380_o;
  wire [1:0] n7382_o;
  wire n7383_o;
  wire [6:0] n7384_o;
  wire n7386_o;
  wire n7387_o;
  wire [2:0] n7388_o;
  wire n7390_o;
  wire n7391_o;
  wire [1:0] n7392_o;
  wire n7394_o;
  wire [2:0] n7395_o;
  wire n7397_o;
  wire n7398_o;
  wire [2:0] n7399_o;
  wire n7401_o;
  wire [1:0] n7402_o;
  wire n7404_o;
  wire n7405_o;
  wire n7406_o;
  wire [2:0] n7407_o;
  wire n7409_o;
  wire n7410_o;
  wire n7411_o;
  wire [1:0] n7412_o;
  wire n7414_o;
  wire n7415_o;
  wire n7418_o;
  wire n7421_o;
  wire n7423_o;
  wire n7426_o;
  wire n7428_o;
  wire n7431_o;
  wire n7434_o;
  wire n7436_o;
  wire n7437_o;
  wire n7438_o;
  wire n7440_o;
  wire n7442_o;
  wire n7444_o;
  wire n7445_o;
  wire [2:0] n7446_o;
  wire n7448_o;
  wire n7449_o;
  wire [1:0] n7450_o;
  wire n7452_o;
  wire [2:0] n7453_o;
  wire n7455_o;
  wire n7456_o;
  wire [2:0] n7457_o;
  wire n7459_o;
  wire [1:0] n7460_o;
  wire n7462_o;
  wire [2:0] n7463_o;
  wire n7465_o;
  wire n7466_o;
  wire n7467_o;
  wire n7468_o;
  wire [4:0] n7469_o;
  wire n7471_o;
  wire [2:0] n7472_o;
  wire n7474_o;
  wire [2:0] n7475_o;
  wire n7477_o;
  wire n7478_o;
  wire [2:0] n7479_o;
  wire n7481_o;
  wire n7484_o;
  wire n7487_o;
  wire n7489_o;
  wire n7492_o;
  wire n7494_o;
  wire n7497_o;
  wire n7500_o;
  wire n7502_o;
  wire n7503_o;
  wire n7504_o;
  wire n7506_o;
  wire n7508_o;
  wire n7510_o;
  wire n7512_o;
  wire n7514_o;
  wire n7516_o;
  wire n7518_o;
  wire n7520_o;
  wire n7522_o;
  wire n7523_o;
  wire n7524_o;
  wire n7525_o;
  wire n7527_o;
  wire [12:0] n7528_o;
  reg n7529_o;
  reg [1:0] n7531_o;
  reg [1:0] n7532_o;
  reg [1:0] n7533_o;
  reg n7534_o;
  reg n7536_o;
  reg n7538_o;
  reg n7540_o;
  reg n7543_o;
  reg n7545_o;
  reg n7547_o;
  reg n7550_o;
  reg n7553_o;
  reg n7556_o;
  reg n7559_o;
  reg n7562_o;
  reg n7565_o;
  reg n7568_o;
  reg n7571_o;
  reg n7574_o;
  reg [1:0] n7576_o;
  reg [5:0] n7577_o;
  reg n7579_o;
  reg n7581_o;
  reg n7584_o;
  reg n7587_o;
  reg n7591_o;
  reg n7594_o;
  reg n7597_o;
  reg n7600_o;
  reg n7606_o;
  reg n7609_o;
  reg n7612_o;
  reg n7615_o;
  reg n7618_o;
  reg n7621_o;
  wire n7623_o;
  reg n7624_o;
  wire [2:0] n7625_o;
  reg [2:0] n7626_o;
  wire n7627_o;
  reg n7628_o;
  wire n7629_o;
  reg n7630_o;
  wire n7631_o;
  reg n7632_o;
  wire n7633_o;
  reg n7634_o;
  wire n7635_o;
  reg n7636_o;
  wire n7637_o;
  reg n7638_o;
  wire n7639_o;
  reg n7640_o;
  reg n7641_o;
  wire n7642_o;
  reg n7643_o;
  wire n7644_o;
  reg n7645_o;
  wire n7646_o;
  wire n7647_o;
  reg n7648_o;
  wire n7649_o;
  wire n7650_o;
  reg n7651_o;
  wire n7652_o;
  reg n7653_o;
  wire n7654_o;
  wire n7655_o;
  wire n7656_o;
  wire n7657_o;
  wire n7658_o;
  reg n7659_o;
  wire n7660_o;
  wire n7661_o;
  wire n7662_o;
  wire n7663_o;
  wire n7664_o;
  reg n7665_o;
  wire n7666_o;
  wire n7667_o;
  reg n7668_o;
  wire n7669_o;
  wire n7670_o;
  reg n7671_o;
  wire n7672_o;
  reg n7673_o;
  wire [1:0] n7674_o;
  wire [1:0] n7675_o;
  reg [1:0] n7676_o;
  wire n7677_o;
  wire n7678_o;
  reg n7679_o;
  wire n7680_o;
  wire n7681_o;
  reg n7682_o;
  wire n7683_o;
  wire n7684_o;
  wire n7685_o;
  reg n7686_o;
  wire n7687_o;
  wire n7688_o;
  reg n7689_o;
  wire [3:0] n7690_o;
  reg [3:0] n7691_o;
  wire n7692_o;
  reg n7693_o;
  wire n7694_o;
  wire [4:0] n7695_o;
  reg [4:0] n7696_o;
  wire n7697_o;
  reg n7698_o;
  wire n7699_o;
  reg n7700_o;
  wire n7701_o;
  reg n7702_o;
  wire n7703_o;
  wire n7704_o;
  reg n7705_o;
  wire n7706_o;
  reg n7707_o;
  wire n7708_o;
  reg n7709_o;
  wire n7710_o;
  reg n7711_o;
  wire n7712_o;
  reg n7713_o;
  wire n7714_o;
  reg n7715_o;
  wire [15:0] n7718_o;
  wire n7719_o;
  wire n7720_o;
  wire [3:0] n7725_o;
  wire n7727_o;
  wire n7731_o;
  wire n7744_o;
  wire n7745_o;
  wire n7746_o;
  wire n7750_o;
  wire n7754_o;
  reg n7756_o;
  wire n7757_o;
  reg n7759_o;
  wire n7760_o;
  reg n7762_o;
  wire n7763_o;
  wire n7764_o;
  reg n7766_o;
  wire n7767_o;
  reg n7769_o;
  wire n7770_o;
  reg n7772_o;
  wire n7773_o;
  wire n7774_o;
  reg n7776_o;
  wire n7777_o;
  wire n7778_o;
  reg n7780_o;
  wire n7781_o;
  reg n7783_o;
  reg n7785_o;
  reg n7787_o;
  reg n7789_o;
  reg n7791_o;
  reg n7793_o;
  reg n7795_o;
  reg n7797_o;
  reg n7799_o;
  reg n7801_o;
  reg n7803_o;
  reg n7805_o;
  reg n7807_o;
  reg [1:0] n7809_o;
  reg n7811_o;
  reg n7813_o;
  reg [1:0] n7815_o;
  reg [1:0] n7817_o;
  reg n7819_o;
  reg n7821_o;
  localparam [88:0] n7822_o = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n7833_o;
  wire [2:0] n7841_o;
  wire n7845_o;
  wire n7847_o;
  wire [31:0] n7852_o;
  wire [6:0] n7854_o;
  wire [1:0] n7857_o;
  wire [5:0] n7858_o;
  reg [6:0] n7859_o;
  wire n7860_o;
  wire n7861_o;
  wire n7862_o;
  wire n7863_o;
  wire [1:0] n7864_o;
  wire n7866_o;
  wire n7867_o;
  wire n7868_o;
  wire n7870_o;
  wire n7871_o;
  wire n7873_o;
  wire n7875_o;
  wire n7877_o;
  wire n7879_o;
  wire n7880_o;
  wire n7882_o;
  wire n7883_o;
  wire n7884_o;
  wire n7885_o;
  wire n7886_o;
  wire n7887_o;
  wire n7888_o;
  wire n7890_o;
  wire n7891_o;
  wire n7892_o;
  wire n7895_o;
  wire [2:0] n7896_o;
  wire n7898_o;
  wire n7900_o;
  wire [1:0] n7904_o;
  wire n7906_o;
  wire n7907_o;
  wire n7908_o;
  wire n7909_o;
  wire [6:0] n7911_o;
  wire n7913_o;
  wire n7914_o;
  wire n7916_o;
  wire n7917_o;
  wire n7918_o;
  wire n7919_o;
  wire n7920_o;
  wire n7921_o;
  wire n7922_o;
  wire n7924_o;
  wire n7926_o;
  wire n7927_o;
  wire n7928_o;
  wire n7929_o;
  wire n7930_o;
  wire n7931_o;
  wire n7932_o;
  wire n7933_o;
  wire n7934_o;
  wire n7935_o;
  wire n7936_o;
  wire n7938_o;
  wire n7939_o;
  wire n7941_o;
  wire n7943_o;
  wire [6:0] n7944_o;
  wire n7945_o;
  wire [6:0] n7947_o;
  wire n7953_o;
  wire n7956_o;
  wire n7959_o;
  wire n7960_o;
  wire n7961_o;
  wire n7963_o;
  wire n7964_o;
  wire n7965_o;
  wire n7967_o;
  wire n7968_o;
  wire n7970_o;
  wire n7971_o;
  wire n7973_o;
  wire n7975_o;
  wire n7976_o;
  wire n7977_o;
  wire n7978_o;
  wire n7979_o;
  wire n7981_o;
  wire [1:0] n7983_o;
  wire n7984_o;
  wire [1:0] n7986_o;
  wire n7989_o;
  wire n7992_o;
  wire n7993_o;
  wire n7994_o;
  wire n7995_o;
  wire n7996_o;
  wire [6:0] n7999_o;
  wire n8001_o;
  wire n8004_o;
  wire n8005_o;
  wire n8008_o;
  wire n8009_o;
  wire n8010_o;
  wire n8011_o;
  wire n8012_o;
  wire n8013_o;
  wire [1:0] n8015_o;
  wire n8017_o;
  wire [6:0] n8020_o;
  wire [1:0] n8021_o;
  wire n8023_o;
  wire [1:0] n8027_o;
  wire n8030_o;
  wire n8032_o;
  wire n8033_o;
  wire n8034_o;
  wire [6:0] n8036_o;
  wire [1:0] n8038_o;
  wire n8040_o;
  wire n8041_o;
  wire n8042_o;
  wire n8043_o;
  wire n8044_o;
  wire [6:0] n8045_o;
  wire n8047_o;
  wire n8050_o;
  wire n8052_o;
  wire n8053_o;
  wire n8054_o;
  wire n8056_o;
  wire [1:0] n8058_o;
  wire n8059_o;
  wire n8061_o;
  wire n8062_o;
  wire n8065_o;
  wire n8066_o;
  wire n8067_o;
  wire n8068_o;
  wire n8069_o;
  wire [1:0] n8073_o;
  wire n8075_o;
  wire n8076_o;
  wire n8077_o;
  wire [6:0] n8079_o;
  wire n8081_o;
  wire n8083_o;
  wire n8084_o;
  wire n8085_o;
  wire n8087_o;
  wire n8088_o;
  wire n8089_o;
  wire n8091_o;
  wire n8092_o;
  wire n8094_o;
  wire n8096_o;
  wire n8097_o;
  wire n8098_o;
  wire n8099_o;
  wire n8101_o;
  wire [1:0] n8103_o;
  wire n8104_o;
  wire [1:0] n8106_o;
  wire n8109_o;
  wire n8112_o;
  wire n8113_o;
  wire n8114_o;
  wire n8115_o;
  wire [6:0] n8118_o;
  wire n8120_o;
  wire n8123_o;
  wire n8124_o;
  wire n8127_o;
  wire n8128_o;
  wire n8129_o;
  wire n8130_o;
  wire n8131_o;
  wire n8132_o;
  wire [1:0] n8134_o;
  wire n8136_o;
  wire [6:0] n8139_o;
  wire [1:0] n8140_o;
  wire n8142_o;
  wire [1:0] n8147_o;
  wire n8148_o;
  wire n8149_o;
  wire n8150_o;
  wire [6:0] n8153_o;
  wire [1:0] n8155_o;
  wire n8156_o;
  wire n8157_o;
  wire n8158_o;
  wire n8159_o;
  wire [6:0] n8160_o;
  wire n8162_o;
  wire n8166_o;
  wire n8169_o;
  wire n8170_o;
  wire n8171_o;
  wire n8173_o;
  wire [1:0] n8175_o;
  wire n8176_o;
  wire n8178_o;
  wire n8180_o;
  wire n8183_o;
  wire n8184_o;
  wire n8185_o;
  wire n8186_o;
  wire n8187_o;
  wire [1:0] n8191_o;
  wire n8192_o;
  wire [6:0] n8195_o;
  wire n8197_o;
  wire n8199_o;
  wire n8202_o;
  wire [6:0] n8204_o;
  wire n8206_o;
  wire n8208_o;
  wire n8209_o;
  wire n8212_o;
  wire n8215_o;
  wire n8217_o;
  wire n8218_o;
  wire n8219_o;
  wire n8221_o;
  wire n8224_o;
  wire [6:0] n8226_o;
  wire n8227_o;
  wire n8230_o;
  wire n8232_o;
  wire n8233_o;
  wire n8235_o;
  wire n8241_o;
  wire n8242_o;
  wire [1:0] n8243_o;
  wire n8245_o;
  wire n8247_o;
  wire n8248_o;
  wire [1:0] n8250_o;
  wire n8253_o;
  wire n8255_o;
  wire n8260_o;
  wire n8262_o;
  wire [1:0] n8264_o;
  wire n8267_o;
  wire n8271_o;
  wire n8272_o;
  wire [1:0] n8274_o;
  wire [6:0] n8276_o;
  wire n8278_o;
  wire n8280_o;
  wire n8281_o;
  wire n8283_o;
  wire n8285_o;
  wire n8287_o;
  wire n8288_o;
  wire [1:0] n8295_o;
  wire n8298_o;
  wire n8299_o;
  wire n8300_o;
  wire n8301_o;
  wire n8302_o;
  wire n8303_o;
  wire n8304_o;
  wire [6:0] n8306_o;
  wire n8308_o;
  wire n8309_o;
  wire n8312_o;
  wire n8318_o;
  wire n8321_o;
  wire n8322_o;
  wire n8324_o;
  wire n8330_o;
  wire n8333_o;
  wire n8334_o;
  wire n8336_o;
  wire [1:0] n8344_o;
  wire n8347_o;
  wire n8349_o;
  wire n8352_o;
  wire n8354_o;
  wire n8355_o;
  wire n8356_o;
  wire n8357_o;
  wire n8358_o;
  wire n8359_o;
  wire n8360_o;
  wire n8361_o;
  wire n8362_o;
  wire n8363_o;
  wire [6:0] n8366_o;
  wire n8368_o;
  wire n8372_o;
  wire n8376_o;
  wire [15:0] n8377_o;
  wire n8379_o;
  wire [2:0] n8380_o;
  wire n8382_o;
  wire n8384_o;
  wire n8386_o;
  wire n8387_o;
  wire n8388_o;
  wire [1:0] n8390_o;
  wire n8391_o;
  wire n8392_o;
  wire [6:0] n8394_o;
  wire n8396_o;
  wire n8397_o;
  wire n8400_o;
  wire n8401_o;
  wire [1:0] n8405_o;
  wire n8406_o;
  wire [1:0] n8408_o;
  wire n8409_o;
  wire n8410_o;
  wire n8411_o;
  wire [6:0] n8413_o;
  wire n8415_o;
  wire [1:0] n8416_o;
  wire n8418_o;
  wire n8420_o;
  wire n8422_o;
  wire [2:0] n8423_o;
  wire n8425_o;
  wire n8427_o;
  wire n8432_o;
  wire [2:0] n8433_o;
  wire n8435_o;
  wire n8437_o;
  wire [1:0] n8439_o;
  wire n8441_o;
  wire [1:0] n8444_o;
  wire n8447_o;
  wire n8449_o;
  wire [2:0] n8450_o;
  wire n8452_o;
  wire n8454_o;
  wire n8457_o;
  wire [2:0] n8458_o;
  wire n8460_o;
  wire n8462_o;
  wire n8465_o;
  wire n8469_o;
  wire n8472_o;
  wire n8475_o;
  wire n8478_o;
  wire n8481_o;
  wire n8484_o;
  wire n8485_o;
  wire n8487_o;
  wire [1:0] n8490_o;
  wire n8491_o;
  wire n8492_o;
  wire [6:0] n8495_o;
  wire n8497_o;
  wire n8498_o;
  wire n8500_o;
  wire n8503_o;
  wire [6:0] n8507_o;
  wire n8509_o;
  wire n8513_o;
  wire n8516_o;
  wire n8519_o;
  wire n8522_o;
  wire n8525_o;
  wire n8526_o;
  wire n8527_o;
  wire n8530_o;
  wire n8531_o;
  wire n8532_o;
  wire n8534_o;
  wire n8536_o;
  wire n8537_o;
  wire n8538_o;
  wire [1:0] n8541_o;
  wire n8543_o;
  wire n8544_o;
  wire [6:0] n8547_o;
  wire n8549_o;
  wire n8551_o;
  wire [3:0] n8552_o;
  wire n8554_o;
  wire [1:0] n8558_o;
  wire [1:0] n8560_o;
  wire n8562_o;
  wire n8563_o;
  wire [6:0] n8566_o;
  wire n8568_o;
  wire n8570_o;
  wire n8572_o;
  wire n8575_o;
  wire [11:0] n8577_o;
  wire n8579_o;
  wire [11:0] n8580_o;
  wire n8582_o;
  wire n8583_o;
  wire [11:0] n8584_o;
  wire n8586_o;
  wire n8587_o;
  wire [11:0] n8588_o;
  wire n8590_o;
  wire n8591_o;
  wire n8592_o;
  wire [11:0] n8593_o;
  wire n8595_o;
  wire [11:0] n8596_o;
  wire n8598_o;
  wire n8599_o;
  wire [11:0] n8600_o;
  wire n8602_o;
  wire n8603_o;
  wire [11:0] n8604_o;
  wire n8606_o;
  wire n8607_o;
  wire n8608_o;
  wire n8609_o;
  wire n8610_o;
  wire n8611_o;
  wire n8613_o;
  wire n8615_o;
  wire n8617_o;
  wire n8618_o;
  wire n8620_o;
  wire n8624_o;
  wire n8626_o;
  wire n8627_o;
  wire n8628_o;
  wire [1:0] n8631_o;
  wire n8633_o;
  wire n8634_o;
  wire n8637_o;
  wire n8638_o;
  wire n8639_o;
  wire n8640_o;
  wire [1:0] n8643_o;
  wire n8645_o;
  wire n8646_o;
  wire n8650_o;
  wire n8651_o;
  wire [1:0] n8654_o;
  wire [1:0] n8656_o;
  wire [1:0] n8657_o;
  wire n8658_o;
  wire n8659_o;
  wire n8660_o;
  wire [6:0] n8662_o;
  wire n8664_o;
  wire n8665_o;
  wire n8666_o;
  wire [1:0] n8669_o;
  wire n8671_o;
  wire n8673_o;
  wire n8674_o;
  wire n8676_o;
  wire [5:0] n8679_o;
  wire n8681_o;
  wire n8684_o;
  wire [6:0] n8687_o;
  wire n8689_o;
  wire n8690_o;
  wire n8691_o;
  wire n8693_o;
  wire n8695_o;
  wire n8696_o;
  wire n8698_o;
  wire n8700_o;
  wire [1:0] n8702_o;
  wire [6:0] n8704_o;
  wire n8706_o;
  wire n8708_o;
  wire n8709_o;
  wire n8710_o;
  wire n8711_o;
  wire n8712_o;
  wire n8714_o;
  wire n8719_o;
  wire n8721_o;
  wire [15:0] n8722_o;
  wire n8724_o;
  wire n8725_o;
  wire n8726_o;
  wire n8728_o;
  wire [15:0] n8729_o;
  wire n8731_o;
  wire n8732_o;
  wire n8735_o;
  wire [6:0] n8737_o;
  wire n8740_o;
  wire n8741_o;
  wire n8743_o;
  wire [5:0] n8746_o;
  wire n8748_o;
  wire n8751_o;
  wire [6:0] n8754_o;
  wire n8756_o;
  wire n8757_o;
  wire n8758_o;
  wire n8759_o;
  wire n8761_o;
  wire n8762_o;
  wire n8763_o;
  wire n8765_o;
  wire [1:0] n8768_o;
  wire n8771_o;
  wire n8772_o;
  wire [6:0] n8774_o;
  wire n8777_o;
  wire n8778_o;
  wire n8781_o;
  wire n8782_o;
  wire n8785_o;
  wire [5:0] n8786_o;
  wire n8788_o;
  wire [5:0] n8789_o;
  wire [5:0] n8791_o;
  wire n8792_o;
  wire n8793_o;
  wire n8795_o;
  wire n8797_o;
  wire [80:0] n8798_o;
  reg n8801_o;
  reg [1:0] n8814_o;
  reg [1:0] n8815_o;
  reg [1:0] n8853_o;
  reg n8856_o;
  reg n8859_o;
  reg n8864_o;
  reg n8866_o;
  reg n8876_o;
  reg n8880_o;
  reg n8894_o;
  reg n8896_o;
  reg n8899_o;
  reg n8902_o;
  reg n8905_o;
  reg n8909_o;
  reg n8913_o;
  reg n8916_o;
  reg n8921_o;
  reg n8923_o;
  reg n8928_o;
  reg n8931_o;
  reg n8937_o;
  reg n8941_o;
  reg n8946_o;
  reg [5:0] n8947_o;
  reg n8951_o;
  reg n8954_o;
  reg n8961_o;
  reg n8963_o;
  reg n8964_o;
  reg n8967_o;
  reg n8969_o;
  reg n8971_o;
  reg n8972_o;
  reg n8973_o;
  reg n8974_o;
  reg n8975_o;
  reg n8976_o;
  reg n8977_o;
  wire n8978_o;
  reg n8979_o;
  reg n8980_o;
  reg n8981_o;
  reg n8982_o;
  reg n8983_o;
  reg n8984_o;
  reg n8985_o;
  reg n8986_o;
  reg n8987_o;
  reg n8988_o;
  reg n8989_o;
  reg n8990_o;
  reg n8991_o;
  reg n8992_o;
  wire n8993_o;
  reg n8994_o;
  wire n8995_o;
  reg n8996_o;
  reg n8997_o;
  wire n8998_o;
  reg n8999_o;
  wire n9000_o;
  reg n9001_o;
  reg n9002_o;
  reg n9003_o;
  reg n9004_o;
  reg n9005_o;
  reg n9006_o;
  wire n9007_o;
  reg n9008_o;
  reg n9009_o;
  reg n9010_o;
  reg n9011_o;
  reg n9012_o;
  reg n9013_o;
  wire n9014_o;
  reg n9015_o;
  wire n9016_o;
  reg n9017_o;
  wire n9018_o;
  wire [1:0] n9020_o;
  wire n9022_o;
  wire [1:0] n9023_o;
  wire [3:0] n9024_o;
  wire n9026_o;
  reg n9027_o;
  wire [1:0] n9028_o;
  wire [1:0] n9029_o;
  reg [6:0] n9070_o;
  wire n9076_o;
  wire n9077_o;
  wire [11:0] n9078_o;
  wire [2:0] n9079_o;
  wire n9081_o;
  wire [2:0] n9082_o;
  wire n9084_o;
  wire [3:0] n9085_o;
  wire n9087_o;
  wire n9089_o;
  wire n9091_o;
  wire n9093_o;
  wire n9095_o;
  wire n9097_o;
  wire [7:0] n9098_o;
  reg [31:0] n9099_o;
  reg [3:0] n9100_o;
  reg [2:0] n9101_o;
  reg [2:0] n9102_o;
  wire [31:0] n9103_o;
  wire [3:0] n9104_o;
  wire [2:0] n9105_o;
  wire [2:0] n9106_o;
  wire [31:0] n9108_o;
  wire [3:0] n9110_o;
  wire [2:0] n9111_o;
  wire [2:0] n9112_o;
  wire [11:0] n9117_o;
  wire [31:0] n9119_o;
  wire n9121_o;
  wire [31:0] n9123_o;
  wire n9125_o;
  wire [3:0] n9127_o;
  wire [31:0] n9129_o;
  wire n9131_o;
  wire n9133_o;
  wire [3:0] n9134_o;
  reg [31:0] n9136_o;
  wire [3:0] n9141_o;
  wire n9143_o;
  wire n9145_o;
  wire n9146_o;
  wire n9147_o;
  wire n9148_o;
  wire n9149_o;
  wire n9150_o;
  wire n9152_o;
  wire n9153_o;
  wire n9154_o;
  wire n9155_o;
  wire n9157_o;
  wire n9158_o;
  wire n9159_o;
  wire n9161_o;
  wire n9162_o;
  wire n9164_o;
  wire n9165_o;
  wire n9166_o;
  wire n9168_o;
  wire n9169_o;
  wire n9171_o;
  wire n9172_o;
  wire n9173_o;
  wire n9175_o;
  wire n9176_o;
  wire n9178_o;
  wire n9179_o;
  wire n9180_o;
  wire n9182_o;
  wire n9183_o;
  wire n9185_o;
  wire n9186_o;
  wire n9187_o;
  wire n9188_o;
  wire n9189_o;
  wire n9190_o;
  wire n9191_o;
  wire n9192_o;
  wire n9193_o;
  wire n9194_o;
  wire n9196_o;
  wire n9197_o;
  wire n9198_o;
  wire n9199_o;
  wire n9200_o;
  wire n9201_o;
  wire n9202_o;
  wire n9203_o;
  wire n9204_o;
  wire n9205_o;
  wire n9207_o;
  wire n9208_o;
  wire n9209_o;
  wire n9210_o;
  wire n9211_o;
  wire n9212_o;
  wire n9213_o;
  wire n9214_o;
  wire n9215_o;
  wire n9216_o;
  wire n9217_o;
  wire n9218_o;
  wire n9219_o;
  wire n9220_o;
  wire n9221_o;
  wire n9222_o;
  wire n9224_o;
  wire n9225_o;
  wire n9226_o;
  wire n9227_o;
  wire n9228_o;
  wire n9229_o;
  wire n9230_o;
  wire n9231_o;
  wire n9232_o;
  wire n9233_o;
  wire n9234_o;
  wire n9235_o;
  wire n9237_o;
  wire [15:0] n9238_o;
  reg n9241_o;
  wire n9246_o;
  wire [15:0] n9247_o;
  wire n9248_o;
  wire n9249_o;
  wire n9250_o;
  wire n9253_o;
  wire n9256_o;
  wire n9259_o;
  wire n9262_o;
  wire n9265_o;
  wire n9268_o;
  wire n9271_o;
  wire n9274_o;
  wire n9277_o;
  wire n9280_o;
  wire n9283_o;
  wire n9286_o;
  wire n9289_o;
  wire n9292_o;
  wire n9295_o;
  wire n9298_o;
  wire [15:0] n9299_o;
  wire n9300_o;
  reg n9301_o;
  wire n9302_o;
  reg n9303_o;
  wire n9304_o;
  reg n9305_o;
  wire n9306_o;
  reg n9307_o;
  wire n9308_o;
  reg n9309_o;
  wire n9310_o;
  reg n9311_o;
  wire n9312_o;
  reg n9313_o;
  wire n9314_o;
  reg n9315_o;
  wire n9316_o;
  reg n9317_o;
  wire n9318_o;
  reg n9319_o;
  wire n9320_o;
  reg n9321_o;
  wire n9322_o;
  reg n9323_o;
  wire n9324_o;
  reg n9325_o;
  wire n9326_o;
  reg n9327_o;
  wire n9328_o;
  reg n9329_o;
  wire n9330_o;
  reg n9331_o;
  wire [15:0] n9332_o;
  wire [15:0] n9333_o;
  wire [15:0] n9334_o;
  wire [3:0] n9342_o;
  wire n9344_o;
  wire [3:0] n9345_o;
  wire n9347_o;
  wire [3:0] n9349_o;
  wire n9351_o;
  wire [3:0] n9352_o;
  wire n9354_o;
  wire n9357_o;
  wire [3:0] n9359_o;
  wire [3:0] n9360_o;
  wire n9362_o;
  wire [3:0] n9363_o;
  wire n9365_o;
  wire [3:0] n9366_o;
  wire [1:0] n9368_o;
  wire n9369_o;
  wire n9370_o;
  wire n9371_o;
  wire n9373_o;
  wire [3:0] n9374_o;
  wire n9376_o;
  wire [3:0] n9377_o;
  wire [1:0] n9378_o;
  wire [1:0] n9380_o;
  localparam [3:0] n9381_o = 4'b0000;
  wire [3:0] n9383_o;
  wire n9385_o;
  wire [1:0] n9387_o;
  wire n9389_o;
  wire n9391_o;
  wire n9392_o;
  wire n9394_o;
  wire n9395_o;
  wire n9396_o;
  wire n9397_o;
  wire n9399_o;
  wire n9400_o;
  wire [1:0] n9401_o;
  wire n9402_o;
  wire n9403_o;
  wire n9404_o;
  wire n9405_o;
  wire n9406_o;
  reg n9409_q;
  wire [3:0] n9410_o;
  reg [3:0] n9411_q;
  wire n9412_o;
  reg n9413_q;
  reg [31:0] n9414_q;
  wire [31:0] n9415_o;
  reg [31:0] n9416_q;
  wire [31:0] n9417_o;
  reg [31:0] n9418_q;
  reg [1:0] n9419_q;
  reg [1:0] n9420_q;
  reg n9421_q;
  reg [15:0] n9422_q;
  reg [15:0] n9423_q;
  wire [15:0] n9424_o;
  reg [15:0] n9425_q;
  reg [31:0] n9426_q;
  reg [31:0] n9427_q;
  reg [15:0] n9428_q;
  wire [3:0] n9430_o;
  reg [3:0] n9431_q;
  wire [31:0] n9432_o;
  wire [3:0] n9435_o;
  reg [3:0] n9436_q;
  wire [3:0] n9437_o;
  reg [3:0] n9438_q;
  wire n9439_o;
  reg n9440_q;
  wire [31:0] n9441_o;
  reg [31:0] n9442_q;
  wire [31:0] n9443_o;
  reg [31:0] n9444_q;
  wire n9445_o;
  reg n9446_q;
  reg [31:0] n9447_q;
  wire [31:0] n9448_o;
  reg [31:0] n9450_q;
  reg n9451_q;
  wire [31:0] n9453_o;
  reg n9454_q;
  reg [15:0] n9455_q;
  reg n9456_q;
  reg n9457_q;
  reg n9458_q;
  reg n9459_q;
  reg n9460_q;
  reg n9461_q;
  reg n9462_q;
  reg [7:0] n9463_q;
  reg n9464_q;
  wire n9465_o;
  reg n9466_q;
  reg [1:0] n9467_q;
  reg [5:0] n9468_q;
  wire n9469_o;
  reg n9470_q;
  wire [3:0] n9471_o;
  reg n9473_q;
  reg n9474_q;
  reg n9475_q;
  reg n9476_q;
  reg n9477_q;
  reg n9478_q;
  reg [7:0] n9479_q;
  reg n9480_q;
  reg n9481_q;
  reg n9482_q;
  reg n9483_q;
  wire [31:0] n9484_o;
  reg [31:0] n9485_q;
  wire [31:0] n9486_o;
  reg [31:0] n9487_q;
  reg [2:0] n9488_q;
  reg [7:0] n9489_q;
  reg n9490_q;
  reg n9491_q;
  reg n9492_q;
  reg n9493_q;
  reg n9494_q;
  wire [31:0] n9495_o;
  wire [7:0] n9496_o;
  reg [7:0] n9497_q;
  reg [5:0] n9498_q;
  reg [3:0] n9499_q;
  reg [5:0] n9500_q;
  reg n9501_q;
  reg n9502_q;
  reg [31:0] n9503_q;
  reg [31:0] n9504_q;
  wire [5:0] n9505_o;
  wire [5:0] n9506_o;
  reg [5:0] n9507_q;
  reg [5:0] n9508_q;
  wire [5:0] n9509_o;
  reg [31:0] n9510_q;
  reg [5:0] n9511_q;
  reg [31:0] n9512_q;
  reg [3:0] n9513_q;
  reg [2:0] n9514_q;
  reg [2:0] n9515_q;
  wire [88:0] n9516_o;
  wire [88:0] n9517_o;
  wire [88:0] n9518_o;
  reg [88:0] n9519_q;
  reg [6:0] n9520_q;
  reg n9521_q;
  reg [1:0] n9522_q;
  wire [2:0] n9523_o;
  wire [31:0] n9525_data; // mem_rd
  wire [31:0] n9526_data; // mem_rd
  assign addr_out = n1035_o;
  assign data_write = n259_o;
  assign nwr = n59_o;
  assign nuds = n70_o;
  assign nlds = n71_o;
  assign busstate = state;
  assign longword = n37_o;
  assign nresetout = n63_o;
  assign fc = n9523_o;
  assign clr_berr = n79_o;
  assign skipFetch = n8801_o;
  assign regin_out = regin;
  assign cacr_out = cacr;
  assign vbr_out = vbr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:148:16  */
  assign use_vbr_stackframe = n9409_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:150:16  */
  assign syncreset = n9411_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:151:16  */
  assign reset = n9413_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:152:16  */
  assign clkena_lw = n75_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:153:16  */
  assign tg68_pc = n9414_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:154:16  */
  assign tmp_tg68_pc = n9416_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:155:16  */
  assign tg68_pc_add = n1136_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:156:16  */
  assign pc_dataa = n1042_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:157:16  */
  assign pc_datab = n1135_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:158:16  */
  assign memaddr = n9418_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:159:16  */
  assign state = n9419_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:160:16  */
  assign datatype = n8814_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:161:16  */
  assign set_datatype = n8815_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:162:16  */
  assign exe_datatype = n9420_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:163:16  */
  assign setstate = n8853_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:164:16  */
  assign setaddrvalue = n8856_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:165:16  */
  assign addrvalue = n9421_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:167:16  */
  assign opcode = n9422_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:168:16  */
  assign exe_opcode = n9423_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:169:16  */
  assign sndopc = n9425_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:171:16  */
  assign exe_pc = n9426_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:172:16  */
  assign last_opc_pc = n9427_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1233:80  */
  assign last_opc_read = n9428_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:175:16  */
  assign reg_qa = n9526_data; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:176:16  */
  assign reg_qb = n9525_data; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:177:16  */
  assign wwrena = n373_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:177:23  */
  assign lwrena = n376_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:178:16  */
  assign bwrena = n379_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:179:16  */
  assign regwrena_now = n8859_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:564:71  */
  assign rf_dest_addr = n421_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:565:73  */
  assign rf_source_addr = n459_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:182:16  */
  assign rf_source_addrd = n9431_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:184:16  */
  assign regin = n9432_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:187:16  */
  assign rdindex_a = n9436_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:188:16  */
  assign rdindex_b = n9438_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:189:16  */
  assign wr_areg = n9440_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:192:16  */
  assign addr = n1034_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:193:16  */
  assign memaddr_reg = n1038_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:194:16  */
  assign memaddr_delta = n1033_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:195:16  */
  assign memaddr_delta_rega = n9442_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:196:16  */
  assign memaddr_delta_regb = n9444_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:197:16  */
  assign use_base = n9446_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:199:16  */
  assign ea_data = n9447_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:200:16  */
  assign op1out = n475_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:201:16  */
  assign op2out = n9448_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:202:16  */
  assign op1outbrief = n800_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:204:16  */
  assign aluout = alu_n23; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:205:16  */
  assign data_write_tmp = n9450_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:206:16  */
  assign data_write_muxin = n222_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:207:16  */
  assign data_write_mux = n231_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:208:16  */
  assign nextpass = n9451_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:209:16  */
  assign setnextpass = n8864_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:210:16  */
  assign setdispbyte = n8866_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:211:16  */
  assign setdisp = n8876_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:212:16  */
  assign regdirectsource = n7536_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:213:16  */
  assign addsub_q = alu_n22; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:214:16  */
  assign briefdata = n836_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:215:16  */
  assign c_out = alu_n21; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:218:16  */
  assign memaddr_a = n9453_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:220:16  */
  assign tg68_pc_brw = n8880_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:221:16  */
  assign tg68_pc_word = n9454_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:222:16  */
  assign getbrief = n7538_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:223:16  */
  assign brief = n9455_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:224:16  */
  assign data_is_source = n7540_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:225:16  */
  assign store_in_tmp = n9456_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:226:16  */
  assign write_back = n7924_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:227:16  */
  assign exec_write_back = n9457_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:228:16  */
  assign setstackaddr = n8894_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:229:16  */
  assign writepc = n8896_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:230:16  */
  assign writepcbig = n9458_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:231:16  */
  assign set_writepcbig = n8899_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:232:16  */
  assign writepcnext = n9459_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:233:16  */
  assign setopcode = n1172_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:234:16  */
  assign decodeopc = n9460_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:235:16  */
  assign execopc = n9461_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:236:16  */
  assign execopc_alu = n41_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:237:16  */
  assign setexecopc = n1197_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:238:16  */
  assign endopc = n9462_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:239:16  */
  assign setendopc = n1176_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:833:98  */
  assign flags = alu_n20; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:241:16  */
  assign flagssr = n9463_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:242:16  */
  assign srin = n1746_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:243:16  */
  assign exec_direct = n9464_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:244:16  */
  assign exec_tas = n9466_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:245:16  */
  assign set_exec_tas = n7550_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:247:16  */
  assign exe_condition = n9241_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:248:16  */
  assign ea_only = n7553_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:249:16  */
  assign source_areg = n8902_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:250:16  */
  assign source_lowbits = n7926_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:251:16  */
  assign source_ldrlbits = n8905_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:252:16  */
  assign source_ldrmbits = n8909_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:253:16  */
  assign source_2ndhbits = n7562_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:254:16  */
  assign source_2ndmbits = n8913_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:255:16  */
  assign source_2ndlbits = n8916_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:256:16  */
  assign dest_areg = n8921_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:257:16  */
  assign dest_ldrareg = n8923_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:258:16  */
  assign dest_ldrhbits = n8928_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:259:16  */
  assign dest_ldrlbits = n8931_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:260:16  */
  assign dest_2ndhbits = n8937_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:261:16  */
  assign dest_2ndlbits = n8941_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:262:16  */
  assign dest_hbits = n8946_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:263:16  */
  assign rot_bits = n9467_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:264:16  */
  assign set_rot_bits = n7576_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:265:16  */
  assign rot_cnt = n9468_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:266:16  */
  assign set_rot_cnt = n8947_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:267:16  */
  assign movem_actiond = n9470_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:268:16  */
  assign movem_regaddr = n9471_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:269:16  */
  assign movem_mux = n9383_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:270:16  */
  assign movem_presub = n7579_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:271:16  */
  assign movem_run = n9385_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:273:16  */
  assign set_direct_data = n8951_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:274:16  */
  assign use_direct_data = n9473_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:275:16  */
  assign direct_data = n9474_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:277:16  */
  assign set_v_flag = alu_n19; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:278:16  */
  assign set_vectoraddr = n8954_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:279:16  */
  assign writesr = n8961_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:280:16  */
  assign trap_berr = n9475_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:281:16  */
  assign trap_illegal = n8963_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:282:16  */
  assign trap_addr_error = 1'b0; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:283:16  */
  assign trap_priv = n7587_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:284:16  */
  assign trap_trace = n9476_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:285:16  */
  assign trap_1010 = n7591_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:286:16  */
  assign trap_1111 = n7594_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:287:16  */
  assign trap_trap = n7597_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:288:16  */
  assign trap_trapv = n7600_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:289:16  */
  assign trap_interrupt = n9477_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:290:16  */
  assign trapmake = n8964_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:291:16  */
  assign trapd = n9478_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:833:79  */
  assign trap_sr = n9479_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:293:16  */
  assign make_trace = n9480_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:294:16  */
  assign make_berr = n9481_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:295:16  */
  assign usestackframe2 = n9482_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:297:16  */
  assign set_stop = n7609_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:298:16  */
  assign stop = n9483_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:299:16  */
  assign trap_vector = n9485_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:300:16  */
  assign trap_vector_vbr = n878_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:301:16  */
  assign usp = n9487_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:306:16  */
  assign ipl_nr = n1199_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:307:16  */
  assign ripl_nr = n9488_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:308:16  */
  assign ipl_vec = n9489_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:309:16  */
  assign interrupt = n9490_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:310:16  */
  assign setinterrupt = n1179_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:311:16  */
  assign svmode = n9491_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:312:16  */
  assign presvmode = n9492_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:313:16  */
  assign suppress_base = n9493_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:314:16  */
  assign set_suppress_base = n8967_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:315:16  */
  assign set_z_error = n8969_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:316:16  */
  assign z_error = n9494_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:317:16  */
  assign ea_build_now = n7890_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:318:16  */
  assign build_logical = n7615_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:319:16  */
  assign build_bcd = n7618_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:321:16  */
  assign data_read = n9495_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:322:16  */
  assign bf_ext_in = n9497_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:323:16  */
  assign bf_ext_out = alu_n17; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:325:16  */
  assign long_start = n215_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:326:16  */
  assign long_start_alu = n39_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:327:16  */
  assign non_aligned = n53_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:328:16  */
  assign check_aligned = n7621_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:329:16  */
  assign long_done = n217_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:330:16  */
  assign memmask = n9498_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:331:16  */
  assign set_memmask = n1730_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:332:16  */
  assign memread = n9499_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:333:16  */
  assign wbmemmask = n9500_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:334:16  */
  assign memmaskmux = n66_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:335:16  */
  assign oddout = n9501_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:336:16  */
  assign set_oddout = n1655_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:337:16  */
  assign pcbase = n9502_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:338:16  */
  assign set_pcbase = n2119_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:340:16  */
  assign last_data_read = n9503_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:341:16  */
  assign last_data_in = n9504_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:343:16  */
  assign bf_offset = n9505_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:344:16  */
  assign bf_width = n9506_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:345:16  */
  assign bf_bhits = n1653_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:346:16  */
  assign bf_shift = n1710_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:347:16  */
  assign alu_width = n9507_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:348:16  */
  assign alu_bf_shift = n9508_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:349:16  */
  assign bf_loffset = n9509_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:350:16  */
  assign bf_full_offset = n1643_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:351:16  */
  assign alu_bf_ffo_offset = n9510_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:352:16  */
  assign alu_bf_loffset = n9511_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:354:16  */
  assign movec_data = n9136_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:355:16  */
  assign vbr = n9512_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:356:16  */
  assign cacr = n9513_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:357:16  */
  assign dfc = n9514_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:358:16  */
  assign sfc = n9515_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:361:16  */
  assign set = n9516_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:362:16  */
  assign set_exec = n9517_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:363:16  */
  assign exec = n9519_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:365:16  */
  assign micro_state = n9520_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:366:16  */
  assign next_micro_state = n9070_o; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:405:49  */
  assign n15_o = last_data_read[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:406:39  */
  assign n16_o = data_read[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:410:31  */
  assign alu_n17 = alu_bf_ext_out; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:414:45  */
  assign n18_o = alu_bf_loffset[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:416:31  */
  assign alu_n19 = alu_set_v_flag; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:417:26  */
  assign alu_n20 = alu_flags; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:418:26  */
  assign alu_n21 = alu_c_out; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:419:29  */
  assign alu_n22 = alu_addsub_q; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:420:27  */
  assign alu_n23 = alu_aluout; // (signal)
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:372:1  */
  tg68k_alu_2_1_2_1 alu (
    .clk(clk),
    .reset(reset),
    .clkena_lw(clkena_lw),
    .cpu(cpu),
    .execopc(execopc_alu),
    .decodeopc(decodeopc),
    .exe_condition(exe_condition),
    .exec_tas(exec_tas),
    .long_start(long_start_alu),
    .non_aligned(non_aligned),
    .check_aligned(check_aligned),
    .movem_presub(movem_presub),
    .set_stop(set_stop),
    .z_error(z_error),
    .rot_bits(rot_bits),
    .exec(exec),
    .op1out(op1out),
    .op2out(op2out),
    .reg_qa(reg_qa),
    .reg_qb(reg_qb),
    .opcode(opcode),
    .exe_opcode(exe_opcode),
    .exe_datatype(exe_datatype),
    .sndopc(sndopc),
    .last_data_read(n15_o),
    .data_read(n16_o),
    .flagssr(flagssr),
    .micro_state(micro_state),
    .bf_ext_in(bf_ext_in),
    .bf_shift(alu_bf_shift),
    .bf_width(alu_width),
    .bf_ffo_offset(alu_bf_ffo_offset),
    .bf_loffset(n18_o),
    .bf_ext_out(alu_bf_ext_out),
    .set_v_flag(alu_set_v_flag),
    .flags(alu_flags),
    .c_out(alu_c_out),
    .addsub_q(alu_addsub_q),
    .aluout(alu_aluout));
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:424:35  */
  assign n36_o = memmaskmux[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:424:21  */
  assign n37_o = ~n36_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:426:48  */
  assign n38_o = memmaskmux[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:426:34  */
  assign n39_o = ~n38_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:427:39  */
  assign n40_o = exec[84];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:427:32  */
  assign n41_o = execopc | n40_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:431:31  */
  assign n44_o = memmaskmux[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:431:44  */
  assign n46_o = n44_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:431:66  */
  assign n47_o = memmaskmux[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:431:79  */
  assign n49_o = n47_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:431:52  */
  assign n50_o = n46_o | n49_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:431:17  */
  assign n53_o = n50_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:441:30  */
  assign n58_o = state == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:441:20  */
  assign n59_o = n58_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:443:35  */
  assign n62_o = exec[74];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:443:26  */
  assign n63_o = n62_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:447:40  */
  assign n65_o = addr[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:447:31  */
  assign n66_o = n65_o ? memmask : n69_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:447:62  */
  assign n67_o = memmask[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:447:75  */
  assign n69_o = {n67_o, 1'b1};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:448:27  */
  assign n70_o = memmaskmux[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:449:27  */
  assign n71_o = memmaskmux[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:450:59  */
  assign n73_o = memmaskmux[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:450:45  */
  assign n74_o = clkena_in & n73_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:450:26  */
  assign n75_o = n74_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:451:44  */
  assign n78_o = setopcode & trap_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:451:25  */
  assign n79_o = n78_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:455:26  */
  assign n83_o = ~nreset;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:460:55  */
  assign n85_o = syncreset[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:460:67  */
  assign n87_o = {n85_o, 1'b1};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:461:55  */
  assign n88_o = syncreset[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:461:42  */
  assign n89_o = ~n88_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:465:52  */
  assign n99_o = cpu[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:465:60  */
  assign n101_o = n99_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:465:45  */
  assign n103_o = 1'b0 | n101_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:465:25  */
  assign n106_o = n103_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:475:30  */
  assign n111_o = memmaskmux[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:475:33  */
  assign n112_o = ~n111_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:476:50  */
  assign n113_o = last_data_in[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:476:63  */
  assign n114_o = {n113_o, data_in};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:478:50  */
  assign n115_o = last_data_in[23:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:478:71  */
  assign n116_o = data_in[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:478:63  */
  assign n117_o = {n115_o, n116_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:480:27  */
  assign n119_o = memread[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:480:46  */
  assign n120_o = memread[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:480:58  */
  assign n122_o = n120_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:480:78  */
  assign n123_o = memmaskmux[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:480:64  */
  assign n124_o = n122_o & n123_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:480:35  */
  assign n125_o = n119_o | n124_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n126_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n127_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n128_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n129_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n130_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n131_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n132_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n133_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n134_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n135_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n136_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n137_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n138_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n139_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n140_o = data_read[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:481:70  */
  assign n141_o = data_read[15];
  assign n142_o = {n126_o, n127_o, n128_o, n129_o};
  assign n143_o = {n130_o, n131_o, n132_o, n133_o};
  assign n144_o = {n134_o, n135_o, n136_o, n137_o};
  assign n145_o = {n138_o, n139_o, n140_o, n141_o};
  assign n146_o = {n142_o, n143_o, n144_o, n145_o};
  assign n147_o = n114_o[31:16];
  assign n148_o = n117_o[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:475:17  */
  assign n149_o = n112_o ? n147_o : n148_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:480:17  */
  assign n150_o = n125_o ? n146_o : n149_o;
  assign n151_o = n114_o[15:0];
  assign n152_o = n117_o[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:475:17  */
  assign n153_o = n112_o ? n151_o : n152_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:485:51  */
  assign n156_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:485:42  */
  assign n157_o = clkena_lw & n156_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:486:46  */
  assign n158_o = memmaskmux[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:486:49  */
  assign n159_o = ~n158_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:487:66  */
  assign n160_o = last_data_in[23:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:489:66  */
  assign n161_o = last_data_in[31:24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:486:33  */
  assign n162_o = n159_o ? n160_o : n161_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:495:41  */
  assign n165_o = state == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:495:54  */
  assign n166_o = exec[38];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:495:47  */
  assign n167_o = n165_o | n166_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:497:49  */
  assign n168_o = state[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:497:52  */
  assign n169_o = ~n168_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:497:68  */
  assign n170_o = memmask[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:497:71  */
  assign n171_o = ~n170_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:497:57  */
  assign n172_o = n169_o & n171_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:499:52  */
  assign n173_o = state[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:499:55  */
  assign n174_o = ~n173_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:499:70  */
  assign n175_o = memread[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:499:60  */
  assign n176_o = n174_o | n175_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n177_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n178_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n179_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n180_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n181_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n182_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n183_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n184_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n185_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n186_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n187_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n188_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n189_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n190_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n191_o = data_in[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:500:97  */
  assign n192_o = data_in[15];
  assign n193_o = {n177_o, n178_o, n179_o, n180_o};
  assign n194_o = {n181_o, n182_o, n183_o, n184_o};
  assign n195_o = {n185_o, n186_o, n187_o, n188_o};
  assign n196_o = {n189_o, n190_o, n191_o, n192_o};
  assign n197_o = {n193_o, n194_o, n195_o, n196_o};
  assign n198_o = data_read[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:499:41  */
  assign n199_o = n176_o ? n197_o : n198_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:497:41  */
  assign n200_o = n172_o ? last_opc_read : n199_o;
  assign n201_o = data_read[15:0];
  assign n202_o = {n200_o, n201_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:494:25  */
  assign n203_o = n206_o ? n202_o : last_data_read;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:503:61  */
  assign n204_o = last_data_in[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:503:74  */
  assign n205_o = {n204_o, data_in};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:494:25  */
  assign n206_o = clkena_in & n167_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:494:25  */
  assign n207_o = clkena_in ? n205_o : last_data_in;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:492:25  */
  assign n209_o = reset ? 32'b00000000000000000000000000000000 : n203_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:492:25  */
  assign n210_o = reset ? last_data_in : n207_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:507:65  */
  assign n214_o = memmask[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:507:54  */
  assign n215_o = ~n214_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:508:64  */
  assign n216_o = memread[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:508:53  */
  assign n217_o = ~n216_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:514:24  */
  assign n221_o = exec[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:514:17  */
  assign n222_o = n221_o ? reg_qb : data_write_tmp;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:527:39  */
  assign n223_o = addr[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:527:34  */
  assign n224_o = oddout == n223_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:528:61  */
  assign n226_o = {8'bX, bf_ext_out};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:528:72  */
  assign n227_o = {n226_o, data_write_muxin};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:530:61  */
  assign n228_o = {bf_ext_out, data_write_muxin};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:530:78  */
  assign n230_o = {n228_o, 8'bX};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:527:25  */
  assign n231_o = n224_o ? n227_o : n230_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:534:30  */
  assign n232_o = memmaskmux[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:534:33  */
  assign n233_o = ~n232_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:535:53  */
  assign n234_o = data_write_mux[47:32];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:536:33  */
  assign n235_o = memmaskmux[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:536:36  */
  assign n236_o = ~n235_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:537:53  */
  assign n237_o = data_write_mux[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:540:38  */
  assign n238_o = memmaskmux[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:540:51  */
  assign n240_o = n238_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:541:61  */
  assign n241_o = data_write_mux[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:541:90  */
  assign n242_o = data_write_mux[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:541:74  */
  assign n243_o = {n241_o, n242_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:542:41  */
  assign n244_o = memmaskmux[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:542:54  */
  assign n246_o = n244_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:543:61  */
  assign n247_o = data_write_mux[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:543:91  */
  assign n248_o = data_write_mux[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:543:75  */
  assign n249_o = {n247_o, n248_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:545:61  */
  assign n250_o = data_write_mux[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:542:25  */
  assign n251_o = n246_o ? n249_o : n250_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:540:25  */
  assign n252_o = n240_o ? n243_o : n251_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:536:17  */
  assign n253_o = n236_o ? n237_o : n252_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:534:17  */
  assign n254_o = n233_o ? n234_o : n253_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:548:24  */
  assign n255_o = exec[72];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:549:53  */
  assign n256_o = data_write_tmp[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:549:83  */
  assign n257_o = data_write_tmp[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:549:67  */
  assign n258_o = {n256_o, n257_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:548:17  */
  assign n259_o = n255_o ? n258_o : n254_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:563:56  */
  assign n272_o = rf_dest_addr[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:570:40  */
  assign n280_o = exec[65];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:561:21  */
  assign n283_o = clkena_lw & wwrena;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:561:21  */
  assign n287_o = clkena_lw & n280_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:583:24  */
  assign n297_o = exec[30];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:585:27  */
  assign n298_o = exec[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:585:44  */
  assign n299_o = n298_o & ea_only;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:587:27  */
  assign n300_o = exec[66];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:589:27  */
  assign n301_o = exec[32];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:594:53  */
  assign n306_o = reg_qa[15:8];
  assign n307_o = memaddr[15:8];
  assign n308_o = memaddr_a[15:8];
  assign n309_o = usp[15:8];
  assign n310_o = movec_data[15:8];
  assign n311_o = aluout[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:589:17  */
  assign n312_o = n301_o ? n310_o : n311_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:587:17  */
  assign n313_o = n300_o ? n309_o : n312_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:585:17  */
  assign n314_o = n299_o ? n308_o : n313_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:583:17  */
  assign n315_o = n297_o ? n307_o : n314_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:593:17  */
  assign n316_o = bwrena ? n306_o : n315_o;
  assign n317_o = memaddr[31:16];
  assign n318_o = memaddr_a[31:16];
  assign n319_o = usp[31:16];
  assign n320_o = movec_data[31:16];
  assign n321_o = aluout[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:589:17  */
  assign n322_o = n301_o ? n320_o : n321_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:587:17  */
  assign n323_o = n300_o ? n319_o : n322_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:585:17  */
  assign n324_o = n299_o ? n318_o : n323_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:583:17  */
  assign n325_o = n297_o ? n317_o : n324_o;
  assign n326_o = memaddr[7:0];
  assign n327_o = memaddr_a[7:0];
  assign n328_o = usp[7:0];
  assign n329_o = movec_data[7:0];
  assign n330_o = aluout[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:589:17  */
  assign n331_o = n301_o ? n329_o : n330_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:587:17  */
  assign n332_o = n300_o ? n328_o : n331_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:585:17  */
  assign n333_o = n299_o ? n327_o : n332_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:583:17  */
  assign n334_o = n297_o ? n326_o : n333_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:596:26  */
  assign n335_o = ~lwrena;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:597:54  */
  assign n336_o = reg_qa[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:596:17  */
  assign n337_o = n335_o ? n336_o : n325_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:24  */
  assign n338_o = exec[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:44  */
  assign n339_o = exec[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:37  */
  assign n340_o = n338_o | n339_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:65  */
  assign n341_o = exec[41];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:58  */
  assign n342_o = n340_o | n341_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:608:27  */
  assign n343_o = exec[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:611:33  */
  assign n345_o = exe_datatype == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:614:56  */
  assign n346_o = wr_areg | movem_actiond;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:614:41  */
  assign n349_o = n346_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:613:33  */
  assign n351_o = exe_datatype == 2'b01;
  assign n352_o = {n351_o, n345_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n352_o)
      2'b10: n355_o = n349_o;
      2'b01: n355_o = 1'b0;
      default: n355_o = 1'b1;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n352_o)
      2'b10: n358_o = 1'b0;
      2'b01: n358_o = 1'b1;
      default: n358_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:608:17  */
  assign n361_o = n343_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:608:17  */
  assign n363_o = n343_o ? n355_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:608:17  */
  assign n365_o = n343_o ? n358_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:606:17  */
  assign n367_o = regwrena_now ? 1'b1 : n361_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:606:17  */
  assign n369_o = regwrena_now ? 1'b0 : n363_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:606:17  */
  assign n371_o = regwrena_now ? 1'b0 : n365_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:17  */
  assign n373_o = n342_o ? 1'b1 : n367_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:17  */
  assign n376_o = n342_o ? 1'b1 : n369_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:603:17  */
  assign n379_o = n342_o ? 1'b0 : n371_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:628:24  */
  assign n384_o = exec[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:630:26  */
  assign n385_o = set[70];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:631:46  */
  assign n386_o = brief[15:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:632:26  */
  assign n387_o = set[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:634:59  */
  assign n388_o = sndopc[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:634:52  */
  assign n390_o = {1'b0, n388_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:639:60  */
  assign n391_o = sndopc[14:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:639:53  */
  assign n392_o = {dest_ldrareg, n391_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:641:55  */
  assign n393_o = last_data_read[15:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:643:59  */
  assign n394_o = last_data_read[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:643:44  */
  assign n396_o = {1'b0, n394_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:645:51  */
  assign n397_o = sndopc[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:645:44  */
  assign n399_o = {1'b0, n397_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:649:57  */
  assign n400_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:649:50  */
  assign n401_o = {dest_areg, n400_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:651:34  */
  assign n402_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:651:46  */
  assign n404_o = n402_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:651:53  */
  assign n405_o = n404_o | data_is_source;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:652:65  */
  assign n406_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:652:58  */
  assign n407_o = {dest_areg, n406_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:654:59  */
  assign n408_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:654:52  */
  assign n410_o = {1'b1, n408_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:651:25  */
  assign n411_o = n405_o ? n407_o : n410_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:648:17  */
  assign n412_o = dest_hbits ? n401_o : n411_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:646:17  */
  assign n414_o = setstackaddr ? 4'b1111 : n412_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:644:17  */
  assign n415_o = dest_2ndlbits ? n399_o : n414_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:642:17  */
  assign n416_o = dest_ldrlbits ? n396_o : n415_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:640:17  */
  assign n417_o = dest_ldrhbits ? n393_o : n416_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:638:17  */
  assign n418_o = dest_2ndhbits ? n392_o : n417_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:632:17  */
  assign n419_o = n387_o ? n390_o : n418_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:630:17  */
  assign n420_o = n385_o ? n386_o : n419_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:628:17  */
  assign n421_o = n384_o ? rf_source_addrd : n420_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:664:24  */
  assign n425_o = exec[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:664:49  */
  assign n426_o = set[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:664:43  */
  assign n427_o = n425_o | n426_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:666:65  */
  assign n429_o = movem_regaddr ^ 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:665:25  */
  assign n430_o = movem_presub ? n429_o : movem_regaddr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:671:53  */
  assign n431_o = sndopc[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:671:46  */
  assign n433_o = {1'b0, n431_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:673:53  */
  assign n434_o = sndopc[14:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:673:46  */
  assign n436_o = {1'b0, n434_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:675:53  */
  assign n437_o = sndopc[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:675:46  */
  assign n439_o = {1'b0, n437_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:677:61  */
  assign n440_o = last_data_read[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:677:46  */
  assign n442_o = {1'b0, n440_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:679:61  */
  assign n443_o = last_data_read[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:679:46  */
  assign n445_o = {1'b0, n443_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:681:61  */
  assign n446_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:681:54  */
  assign n447_o = {source_areg, n446_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:682:27  */
  assign n448_o = exec[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:685:61  */
  assign n449_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:685:54  */
  assign n450_o = {source_areg, n449_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:682:17  */
  assign n452_o = n448_o ? 4'b1111 : n450_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:680:17  */
  assign n453_o = source_lowbits ? n447_o : n452_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:678:17  */
  assign n454_o = source_ldrmbits ? n445_o : n453_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:676:17  */
  assign n455_o = source_ldrlbits ? n442_o : n454_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:674:17  */
  assign n456_o = source_2ndmbits ? n439_o : n455_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:672:17  */
  assign n457_o = source_2ndhbits ? n436_o : n456_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:670:17  */
  assign n458_o = source_2ndlbits ? n433_o : n457_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:664:17  */
  assign n459_o = n427_o ? n430_o : n458_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:695:24  */
  assign n463_o = exec[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:697:27  */
  assign n464_o = exec[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:697:45  */
  assign n465_o = n464_o & store_in_tmp;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:699:27  */
  assign n466_o = exec[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:699:59  */
  assign n467_o = memmaskmux[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:699:62  */
  assign n468_o = ~n467_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:699:46  */
  assign n469_o = n466_o | n468_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:699:74  */
  assign n470_o = exec[39];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:699:67  */
  assign n471_o = n469_o | n470_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:699:17  */
  assign n472_o = n471_o ? addr : reg_qa;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:697:17  */
  assign n473_o = n465_o ? ea_data : n472_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:695:17  */
  assign n475_o = n463_o ? 32'b00000000000000000000000000000000 : n473_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:710:46  */
  assign n479_o = reg_qb[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n480_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n481_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n482_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n483_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n484_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n485_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n486_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n487_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n488_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n489_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n490_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n491_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n492_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n493_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n494_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:711:58  */
  assign n495_o = op2out[15];
  assign n496_o = {n480_o, n481_o, n482_o, n483_o};
  assign n497_o = {n484_o, n485_o, n486_o, n487_o};
  assign n498_o = {n488_o, n489_o, n490_o, n491_o};
  assign n499_o = {n492_o, n493_o, n494_o, n495_o};
  assign n500_o = {n496_o, n497_o, n498_o, n499_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:712:24  */
  assign n501_o = exec[53];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:51  */
  assign n503_o = exec[61];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:61  */
  assign n504_o = n503_o & execopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:43  */
  assign n505_o = use_direct_data | n504_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:85  */
  assign n506_o = exec[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:78  */
  assign n507_o = n505_o | n506_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:28  */
  assign n508_o = exec[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:41  */
  assign n509_o = ~n508_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:46  */
  assign n510_o = n509_o & store_in_tmp;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:75  */
  assign n511_o = exec[27];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:68  */
  assign n512_o = n510_o | n511_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:718:27  */
  assign n513_o = exec[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:719:57  */
  assign n514_o = exe_opcode[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n515_o = exe_opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n516_o = exe_opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n517_o = exe_opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n518_o = exe_opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n519_o = exe_opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n520_o = exe_opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n521_o = exe_opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:720:69  */
  assign n522_o = exe_opcode[7];
  assign n523_o = {n515_o, n516_o, n517_o, n518_o};
  assign n524_o = {n519_o, n520_o, n521_o, n522_o};
  assign n525_o = {n523_o, n524_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:721:27  */
  assign n526_o = exec[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:722:57  */
  assign n527_o = exe_opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:723:38  */
  assign n528_o = exe_opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:723:51  */
  assign n530_o = n528_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:723:25  */
  assign n533_o = n530_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:729:35  */
  assign n536_o = exe_datatype == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:729:49  */
  assign n537_o = exec[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:729:57  */
  assign n538_o = ~n537_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:729:41  */
  assign n539_o = n536_o & n538_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:730:55  */
  assign n540_o = reg_qb[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:729:17  */
  assign n541_o = n539_o ? n540_o : n500_o;
  assign n542_o = {12'b000000000000, n533_o, n527_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:721:17  */
  assign n543_o = n526_o ? n542_o : n479_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:721:17  */
  assign n544_o = n526_o ? n500_o : n541_o;
  assign n545_o = {n544_o, n543_o};
  assign n546_o = {n525_o, n514_o};
  assign n547_o = n545_o[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:718:17  */
  assign n548_o = n513_o ? n546_o : n547_o;
  assign n549_o = n545_o[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:718:17  */
  assign n550_o = n513_o ? n500_o : n549_o;
  assign n551_o = {n550_o, n548_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:17  */
  assign n552_o = n512_o ? ea_data : n551_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:17  */
  assign n553_o = n507_o ? data_write_tmp : n552_o;
  assign n556_o = n553_o[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:712:17  */
  assign n557_o = n501_o ? n500_o : n556_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:732:24  */
  assign n558_o = exec[88];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n559_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n560_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n561_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n562_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n563_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n564_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n565_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n566_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n567_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n568_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n569_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n570_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n571_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n572_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n573_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n574_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n575_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n576_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n577_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n578_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n579_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n580_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n581_o = op2out[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:733:65  */
  assign n582_o = op2out[7];
  assign n583_o = {n559_o, n560_o, n561_o, n562_o};
  assign n584_o = {n563_o, n564_o, n565_o, n566_o};
  assign n585_o = {n567_o, n568_o, n569_o, n570_o};
  assign n586_o = {n571_o, n572_o, n573_o, n574_o};
  assign n587_o = {n575_o, n576_o, n577_o, n578_o};
  assign n588_o = {n579_o, n580_o, n581_o, n582_o};
  assign n589_o = {n583_o, n584_o, n585_o, n586_o};
  assign n590_o = {n587_o, n588_o};
  assign n591_o = {n589_o, n590_o};
  assign n592_o = n502_o[15:8];
  assign n593_o = data_write_tmp[15:8];
  assign n594_o = ea_data[15:8];
  assign n595_o = n551_o[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:17  */
  assign n596_o = n512_o ? n594_o : n595_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:17  */
  assign n597_o = n507_o ? n593_o : n596_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:712:17  */
  assign n598_o = n501_o ? n592_o : n597_o;
  assign n599_o = {n557_o, n598_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:732:17  */
  assign n600_o = n558_o ? n591_o : n599_o;
  assign n601_o = n502_o[7:0];
  assign n602_o = data_write_tmp[7:0];
  assign n603_o = ea_data[7:0];
  assign n604_o = n551_o[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:716:17  */
  assign n605_o = n512_o ? n603_o : n604_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:714:17  */
  assign n606_o = n507_o ? n602_o : n605_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:712:17  */
  assign n607_o = n501_o ? n601_o : n606_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:753:40  */
  assign n612_o = exec[82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:753:33  */
  assign n614_o = n612_o ? 1'b1 : use_direct_data;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:759:56  */
  assign n615_o = set[27];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:759:50  */
  assign n616_o = endopc | n615_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:759:33  */
  assign n618_o = n616_o ? 1'b0 : n614_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:756:33  */
  assign n620_o = set_direct_data ? 1'b1 : n618_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:756:33  */
  assign n623_o = set_direct_data ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:762:56  */
  assign n625_o = set_exec[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:769:41  */
  assign n627_o = set_z_error ? 1'b1 : z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:772:52  */
  assign n628_o = set_exec[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:772:75  */
  assign n630_o = state == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:772:66  */
  assign n631_o = n628_o & n630_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:772:41  */
  assign n633_o = n631_o ? 1'b1 : n620_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:776:49  */
  assign n635_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:776:62  */
  assign n636_o = exec[80];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:776:55  */
  assign n637_o = n635_o | n636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:776:41  */
  assign n639_o = n637_o ? 1'b1 : store_in_tmp;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:779:69  */
  assign n641_o = state == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:779:60  */
  assign n642_o = direct_data & n641_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:779:41  */
  assign n644_o = n642_o ? 1'b1 : n639_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:764:33  */
  assign n646_o = endopc ? 1'b0 : n644_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:764:33  */
  assign n648_o = endopc ? 1'b0 : writepcnext;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:764:33  */
  assign n649_o = endopc ? n620_o : n633_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:764:33  */
  assign n651_o = endopc ? 1'b0 : n627_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:784:41  */
  assign n653_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:784:55  */
  assign n654_o = exec[79];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:784:69  */
  assign n655_o = ~n654_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:784:47  */
  assign n656_o = n653_o & n655_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:786:43  */
  assign n657_o = exec[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:788:43  */
  assign n658_o = exec[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:788:92  */
  assign n660_o = state == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:788:83  */
  assign n661_o = direct_data & n660_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:788:63  */
  assign n662_o = n658_o | n661_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:788:33  */
  assign n663_o = n662_o ? last_data_read : ea_data;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:786:33  */
  assign n664_o = n657_o ? addr : n663_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:784:33  */
  assign n665_o = n656_o ? data_read : n664_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:794:43  */
  assign n666_o = exec[25];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:797:50  */
  assign n668_o = micro_state == 7'b0110010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:800:66  */
  assign n669_o = trap_trap | trap_trapv;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:800:87  */
  assign n670_o = exec[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:800:80  */
  assign n671_o = n669_o | n670_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:800:98  */
  assign n672_o = n671_o | z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:801:51  */
  assign n674_o = micro_state == 7'b0110011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:807:100  */
  assign n675_o = trap_vector[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:807:87  */
  assign n677_o = {4'b0010, n675_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:809:100  */
  assign n678_o = trap_vector[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:809:87  */
  assign n680_o = {4'b0000, n678_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:810:74  */
  assign n681_o = trap_trap | trap_trapv;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:810:95  */
  assign n682_o = exec[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:810:88  */
  assign n683_o = n681_o | n682_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:810:106  */
  assign n684_o = n683_o | z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:805:41  */
  assign n685_o = usestackframe2 ? n677_o : n680_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:805:41  */
  assign n686_o = usestackframe2 ? n648_o : n684_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:815:43  */
  assign n687_o = exec[64];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:817:43  */
  assign n688_o = exec[61];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:819:43  */
  assign n689_o = exec[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:819:60  */
  assign n690_o = n689_o & ea_only;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:823:65  */
  assign n692_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:823:56  */
  assign n693_o = exec_direct & n692_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:825:49  */
  assign n694_o = exec[37];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:826:94  */
  assign n695_o = data_write_tmp[23:0];
  assign n696_o = data_read[31:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:825:41  */
  assign n697_o = n694_o ? n695_o : n696_o;
  assign n698_o = data_read[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:828:43  */
  assign n699_o = exec[37];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:829:78  */
  assign n700_o = reg_qb[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:833:91  */
  assign n701_o = {trap_sr, flags};
  assign n702_o = op2out[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:832:33  */
  assign n703_o = writesr ? n701_o : n702_o;
  assign n704_o = op2out[31:16];
  assign n705_o = data_write_tmp[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:832:33  */
  assign n706_o = writesr ? n705_o : n704_o;
  assign n707_o = {n706_o, n703_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:830:33  */
  assign n708_o = direct_data ? last_data_read : n707_o;
  assign n709_o = n708_o[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:828:33  */
  assign n710_o = n699_o ? n700_o : n709_o;
  assign n711_o = n708_o[31:16];
  assign n712_o = data_write_tmp[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:828:33  */
  assign n713_o = n699_o ? n712_o : n711_o;
  assign n714_o = {n713_o, n710_o};
  assign n715_o = {n697_o, n698_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:823:33  */
  assign n716_o = n693_o ? n715_o : n714_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:821:33  */
  assign n717_o = execopc ? aluout : n716_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:819:33  */
  assign n718_o = n690_o ? addr : n717_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:817:33  */
  assign n719_o = n688_o ? op1out : n718_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:815:33  */
  assign n720_o = n687_o ? data_write_tmp : n719_o;
  assign n721_o = n720_o[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:801:33  */
  assign n722_o = n674_o ? n685_o : n721_o;
  assign n723_o = n720_o[31:16];
  assign n724_o = data_write_tmp[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:801:33  */
  assign n725_o = n674_o ? n724_o : n723_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:801:33  */
  assign n726_o = n674_o ? n686_o : n648_o;
  assign n727_o = {n725_o, n722_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:797:33  */
  assign n728_o = n668_o ? exe_pc : n727_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:797:33  */
  assign n729_o = n668_o ? n672_o : n726_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:797:33  */
  assign n732_o = n668_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:794:33  */
  assign n733_o = n666_o ? tg68_pc_add : n728_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:794:33  */
  assign n734_o = n666_o ? n648_o : n729_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:794:33  */
  assign n736_o = n666_o ? 1'b0 : n732_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:792:33  */
  assign n737_o = writepc ? tg68_pc : n733_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:792:33  */
  assign n738_o = writepc ? n648_o : n734_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:792:33  */
  assign n740_o = writepc ? 1'b0 : n736_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n742_o = clkena_lw ? n665_o : ea_data;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n743_o = clkena_lw ? n737_o : data_write_tmp;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n744_o = clkena_lw ? n646_o : store_in_tmp;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n745_o = clkena_lw ? n738_o : writepcnext;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n746_o = clkena_lw ? n625_o : exec_direct;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n747_o = clkena_lw ? n649_o : use_direct_data;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n748_o = clkena_lw ? n623_o : direct_data;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n749_o = clkena_lw ? n740_o : usestackframe2;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:750:25  */
  assign n750_o = clkena_lw ? n651_o : z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n751_o = reset ? ea_data : n742_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n752_o = reset ? data_write_tmp : n743_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n754_o = reset ? 1'b0 : n744_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n756_o = reset ? 1'b0 : n745_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n757_o = reset ? exec_direct : n746_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n759_o = reset ? 1'b0 : n747_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n761_o = reset ? 1'b0 : n748_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n762_o = reset ? usestackframe2 : n749_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:744:25  */
  assign n764_o = reset ? 1'b0 : n750_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:846:25  */
  assign n777_o = brief[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:847:46  */
  assign n778_o = op1out[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n779_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n780_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n781_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n782_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n783_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n784_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n785_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n786_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n787_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n788_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n789_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n790_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n791_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n792_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n793_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:849:55  */
  assign n794_o = op1out[15];
  assign n795_o = {n779_o, n780_o, n781_o, n782_o};
  assign n796_o = {n783_o, n784_o, n785_o, n786_o};
  assign n797_o = {n787_o, n788_o, n789_o, n790_o};
  assign n798_o = {n791_o, n792_o, n793_o, n794_o};
  assign n799_o = {n795_o, n796_o, n797_o, n798_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:846:17  */
  assign n800_o = n777_o ? n778_o : n799_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:851:48  */
  assign n801_o = op1out[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:851:41  */
  assign n802_o = {op1outbrief, n801_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:852:42  */
  assign n803_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:852:50  */
  assign n805_o = n803_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:852:35  */
  assign n807_o = 1'b0 | n805_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:853:35  */
  assign n808_o = brief[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:854:77  */
  assign n809_o = op1out[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:854:70  */
  assign n810_o = {op1outbrief, n809_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:854:33  */
  assign n812_o = n808_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:855:70  */
  assign n813_o = op1outbrief[14:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:855:90  */
  assign n814_o = op1out[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:855:83  */
  assign n815_o = {n813_o, n814_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:855:103  */
  assign n817_o = {n815_o, 1'b0};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:855:33  */
  assign n819_o = n808_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:856:70  */
  assign n820_o = op1outbrief[13:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:856:90  */
  assign n821_o = op1out[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:856:83  */
  assign n822_o = {n820_o, n821_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:856:103  */
  assign n824_o = {n822_o, 2'b00};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:856:33  */
  assign n826_o = n808_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:857:70  */
  assign n827_o = op1outbrief[12:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:857:90  */
  assign n828_o = op1out[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:857:83  */
  assign n829_o = {n827_o, n828_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:857:103  */
  assign n831_o = {n829_o, 3'b000};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:857:33  */
  assign n833_o = n808_o == 2'b11;
  assign n834_o = {n833_o, n826_o, n819_o, n812_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:853:25  */
  always @*
    case (n834_o)
      4'b1000: n835_o = n831_o;
      4'b0100: n835_o = n824_o;
      4'b0010: n835_o = n817_o;
      4'b0001: n835_o = n810_o;
      default: n835_o = n802_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:852:17  */
  assign n836_o = n807_o ? n835_o : n802_o;
  assign n843_o = trap_vector[9:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:873:33  */
  assign n844_o = trap_berr ? 10'b0000001000 : n843_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:876:33  */
  assign n846_o = trap_addr_error ? 10'b0000001100 : n844_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:879:33  */
  assign n848_o = trap_illegal ? 10'b0000010000 : n846_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:882:33  */
  assign n850_o = set_z_error ? 10'b0000010100 : n848_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:885:40  */
  assign n851_o = exec[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:885:33  */
  assign n853_o = n851_o ? 10'b0000011000 : n850_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:888:33  */
  assign n855_o = trap_trapv ? 10'b0000011100 : n853_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:891:33  */
  assign n857_o = trap_priv ? 10'b0000100000 : n855_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:894:33  */
  assign n859_o = trap_trace ? 10'b0000100100 : n857_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:897:33  */
  assign n861_o = trap_1010 ? 10'b0000101000 : n859_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:900:33  */
  assign n863_o = trap_1111 ? 10'b0000101100 : n861_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:904:83  */
  assign n864_o = opcode[3:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:904:75  */
  assign n866_o = {4'b0010, n864_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:904:96  */
  assign n868_o = {n866_o, 2'b00};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:903:33  */
  assign n869_o = trap_trap ? n868_o : n863_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:906:55  */
  assign n870_o = trap_interrupt | set_vectoraddr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:907:76  */
  assign n872_o = {ipl_vec, 2'b00};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:906:33  */
  assign n873_o = n870_o ? n872_o : n869_o;
  assign n874_o = {22'b0000000000000000000000, n873_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:912:55  */
  assign n877_o = trap_vector + vbr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:911:17  */
  assign n878_o = use_vbr_stackframe ? n877_o : trap_vector;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:918:60  */
  assign n880_o = memaddr_a[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:918:60  */
  assign n881_o = memaddr_a[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:918:60  */
  assign n882_o = memaddr_a[4];
  assign n883_o = {n880_o, n881_o, n882_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n884_o = memaddr_a[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n885_o = memaddr_a[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n886_o = memaddr_a[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n887_o = memaddr_a[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n888_o = memaddr_a[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n889_o = memaddr_a[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n890_o = memaddr_a[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:919:61  */
  assign n891_o = memaddr_a[7];
  assign n892_o = {n884_o, n885_o, n886_o, n887_o};
  assign n893_o = {n888_o, n889_o, n890_o, n891_o};
  assign n894_o = {n892_o, n893_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n895_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n896_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n897_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n898_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n899_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n900_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n901_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n902_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n903_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n904_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n905_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n906_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n907_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n908_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n909_o = memaddr_a[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:920:62  */
  assign n910_o = memaddr_a[15];
  assign n911_o = {n895_o, n896_o, n897_o, n898_o};
  assign n912_o = {n899_o, n900_o, n901_o, n902_o};
  assign n913_o = {n903_o, n904_o, n905_o, n906_o};
  assign n914_o = {n907_o, n908_o, n909_o, n910_o};
  assign n915_o = {n911_o, n912_o, n913_o, n914_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:922:32  */
  assign n916_o = exec[70];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:923:55  */
  assign n917_o = briefdata + memaddr_delta;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:925:72  */
  assign n918_o = last_data_read[7:0];
  assign n919_o = last_data_read[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:924:25  */
  assign n920_o = setdispbyte ? n918_o : n919_o;
  assign n921_o = last_data_read[31:8];
  assign n922_o = {n915_o, n894_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:924:25  */
  assign n923_o = setdispbyte ? n922_o : n921_o;
  assign n924_o = {n923_o, n920_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:922:25  */
  assign n925_o = n916_o ? n917_o : n924_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:929:26  */
  assign n926_o = set[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:930:31  */
  assign n927_o = set[73];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:932:39  */
  assign n930_o = datatype == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:932:52  */
  assign n931_o = set[50];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:932:60  */
  assign n932_o = ~n931_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:932:45  */
  assign n933_o = n930_o & n932_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:932:25  */
  assign n936_o = n933_o ? 5'b11111 : 5'b11110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:930:25  */
  assign n937_o = n927_o ? 5'b11100 : n936_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:938:53  */
  assign n939_o = {1'b1, ripl_nr};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:938:61  */
  assign n941_o = {n939_o, 1'b0};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:937:17  */
  assign n942_o = interrupt ? n941_o : 5'b00000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:929:17  */
  assign n943_o = n926_o ? n937_o : n942_o;
  assign n944_o = n925_o[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:921:17  */
  assign n945_o = setdisp ? n944_o : n943_o;
  assign n946_o = n925_o[31:5];
  assign n947_o = {n915_o, n894_o, n883_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:921:17  */
  assign n948_o = setdisp ? n946_o : n947_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:943:40  */
  assign n950_o = exec[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:943:66  */
  assign n952_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:943:83  */
  assign n953_o = memread[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:943:72  */
  assign n954_o = n952_o & n953_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:943:57  */
  assign n955_o = n950_o | n954_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:948:46  */
  assign n957_o = memmaskmux[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:948:49  */
  assign n958_o = ~n957_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:948:61  */
  assign n959_o = exec[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:948:54  */
  assign n960_o = n958_o | n959_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:950:42  */
  assign n961_o = set[83];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:952:43  */
  assign n962_o = exec[58];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:954:43  */
  assign n963_o = exec[63];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:954:70  */
  assign n965_o = setstate == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:954:58  */
  assign n966_o = n963_o & n965_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:956:42  */
  assign n967_o = set[45];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:958:47  */
  assign n969_o = setstate == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:960:43  */
  assign n970_o = exec[22];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:967:53  */
  assign n971_o = ~interrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:967:75  */
  assign n972_o = ~suppress_base;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:967:58  */
  assign n973_o = n971_o & n972_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:967:41  */
  assign n976_o = n973_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:963:33  */
  assign n977_o = set_vectoraddr ? trap_vector_vbr : memaddr_a;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:963:33  */
  assign n979_o = set_vectoraddr ? 1'b0 : n976_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:960:33  */
  assign n980_o = n970_o ? ea_data : n977_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:960:33  */
  assign n982_o = n970_o ? memaddr_a : 32'b00000000000000000000000000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:960:33  */
  assign n984_o = n970_o ? 1'b0 : n979_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:958:33  */
  assign n985_o = n969_o ? tg68_pc_add : n980_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:958:33  */
  assign n987_o = n969_o ? 32'b00000000000000000000000000000000 : n982_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:958:33  */
  assign n989_o = n969_o ? 1'b0 : n984_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:956:33  */
  assign n990_o = n967_o ? last_data_read : n985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:956:33  */
  assign n992_o = n967_o ? 32'b00000000000000000000000000000000 : n987_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:956:33  */
  assign n994_o = n967_o ? 1'b0 : n989_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:954:33  */
  assign n995_o = n966_o ? addr : n990_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:954:33  */
  assign n997_o = n966_o ? 32'b00000000000000000000000000000000 : n992_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:954:33  */
  assign n999_o = n966_o ? 1'b0 : n994_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:952:33  */
  assign n1000_o = n962_o ? data_read : n995_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:952:33  */
  assign n1002_o = n962_o ? 32'b00000000000000000000000000000000 : n997_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:952:33  */
  assign n1004_o = n962_o ? 1'b0 : n999_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:950:33  */
  assign n1005_o = n961_o ? tmp_tg68_pc : n1000_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:950:33  */
  assign n1007_o = n961_o ? 32'b00000000000000000000000000000000 : n1002_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:950:33  */
  assign n1009_o = n961_o ? 1'b0 : n1004_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:948:33  */
  assign n1010_o = n960_o ? addsub_q : n1005_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:948:33  */
  assign n1012_o = n960_o ? 32'b00000000000000000000000000000000 : n1007_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:948:33  */
  assign n1015_o = n960_o ? 1'b0 : n1009_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:975:53  */
  assign n1017_o = memread[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:975:73  */
  assign n1018_o = state[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:975:64  */
  assign n1019_o = n1017_o & n1018_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:975:100  */
  assign n1020_o = ~movem_presub;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:975:84  */
  assign n1021_o = n1019_o | n1020_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:942:25  */
  assign n1023_o = clkena_in & n955_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:942:25  */
  assign n1024_o = clkena_in & n1021_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:981:53  */
  assign n1033_o = memaddr_delta_rega + memaddr_delta_regb;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:983:36  */
  assign n1034_o = memaddr_reg + memaddr_delta;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:984:41  */
  assign n1035_o = memaddr_reg + memaddr_delta;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:986:28  */
  assign n1036_o = ~use_base;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:986:17  */
  assign n1038_o = n1036_o ? 32'b00000000000000000000000000000000 : reg_qa;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1001:17  */
  assign n1042_o = tg68_pc_brw ? tmp_tg68_pc : tg68_pc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1006:40  */
  assign n1044_o = pc_datab[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1007:60  */
  assign n1045_o = pc_datab[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1007:60  */
  assign n1046_o = pc_datab[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1007:60  */
  assign n1047_o = pc_datab[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1007:60  */
  assign n1048_o = pc_datab[3];
  assign n1049_o = {n1045_o, n1046_o, n1047_o, n1048_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1050_o = pc_datab[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1051_o = pc_datab[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1052_o = pc_datab[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1053_o = pc_datab[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1054_o = pc_datab[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1055_o = pc_datab[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1056_o = pc_datab[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1008:61  */
  assign n1057_o = pc_datab[7];
  assign n1058_o = {n1050_o, n1051_o, n1052_o, n1053_o};
  assign n1059_o = {n1054_o, n1055_o, n1056_o, n1057_o};
  assign n1060_o = {n1058_o, n1059_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1061_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1062_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1063_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1064_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1065_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1066_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1067_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1068_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1069_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1070_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1071_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1072_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1073_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1074_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1075_o = pc_datab[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1009:62  */
  assign n1076_o = pc_datab[15];
  assign n1077_o = {n1061_o, n1062_o, n1063_o, n1064_o};
  assign n1078_o = {n1065_o, n1066_o, n1067_o, n1068_o};
  assign n1079_o = {n1069_o, n1070_o, n1071_o, n1072_o};
  assign n1080_o = {n1073_o, n1074_o, n1075_o, n1076_o};
  assign n1081_o = {n1077_o, n1078_o, n1079_o, n1080_o};
  assign n1085_o = n1043_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1013:24  */
  assign n1086_o = exec[25];
  assign n1090_o = n1082_o[0];
  assign n1091_o = n1043_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1010:17  */
  assign n1092_o = interrupt ? n1090_o : n1091_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1014:25  */
  assign n1093_o = writepcbig ? 1'b1 : n1092_o;
  assign n1094_o = n1082_o[1];
  assign n1095_o = n1043_o[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1010:17  */
  assign n1096_o = interrupt ? n1094_o : n1095_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1014:25  */
  assign n1097_o = writepcbig ? n1096_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1014:25  */
  assign n1098_o = writepcbig ? 1'b1 : n1044_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:47  */
  assign n1099_o = ~use_vbr_stackframe;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:71  */
  assign n1100_o = trap_trap | trap_trapv;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:96  */
  assign n1101_o = exec[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:89  */
  assign n1102_o = n1100_o | n1101_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:111  */
  assign n1103_o = n1102_o | z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:52  */
  assign n1104_o = n1099_o & n1103_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:128  */
  assign n1105_o = n1104_o | writepcnext;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1020:25  */
  assign n1107_o = n1105_o ? 1'b1 : n1093_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1023:28  */
  assign n1109_o = state == 2'b00;
  assign n1111_o = n1082_o[0];
  assign n1112_o = n1043_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1010:17  */
  assign n1113_o = interrupt ? n1111_o : n1112_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1023:17  */
  assign n1114_o = n1109_o ? 1'b1 : n1113_o;
  assign n1115_o = {n1098_o, n1097_o, n1107_o};
  assign n1116_o = n1115_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1013:17  */
  assign n1117_o = n1086_o ? n1116_o : n1114_o;
  assign n1118_o = n1115_o[2:1];
  assign n1119_o = n1082_o[1];
  assign n1120_o = n1043_o[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1010:17  */
  assign n1121_o = interrupt ? n1119_o : n1120_o;
  assign n1122_o = {n1044_o, n1121_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1013:17  */
  assign n1123_o = n1086_o ? n1118_o : n1122_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1030:63  */
  assign n1127_o = opcode[7:0];
  assign n1128_o = last_data_read[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1027:25  */
  assign n1129_o = tg68_pc_word ? n1128_o : n1127_o;
  assign n1130_o = last_data_read[31:8];
  assign n1131_o = {n1081_o, n1060_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1027:25  */
  assign n1132_o = tg68_pc_word ? n1130_o : n1131_o;
  assign n1133_o = {n1132_o, n1129_o};
  assign n1134_o = {n1081_o, n1060_o, n1049_o, n1123_o, n1117_o, n1085_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1026:17  */
  assign n1135_o = tg68_pc_brw ? n1133_o : n1134_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1034:40  */
  assign n1136_o = pc_dataa + pc_datab;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:28  */
  assign n1138_o = setstate == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:54  */
  assign n1140_o = next_micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:34  */
  assign n1141_o = n1138_o & n1140_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:75  */
  assign n1142_o = ~setnextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:60  */
  assign n1143_o = n1141_o & n1142_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:100  */
  assign n1144_o = ~exec_write_back;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:113  */
  assign n1146_o = state == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:105  */
  assign n1147_o = n1144_o | n1146_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:80  */
  assign n1148_o = n1143_o & n1147_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:135  */
  assign n1150_o = set_rot_cnt == 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:120  */
  assign n1151_o = n1148_o & n1150_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:157  */
  assign n1152_o = set_exec[31];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:165  */
  assign n1153_o = ~n1152_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:145  */
  assign n1154_o = n1151_o & n1153_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:35  */
  assign n1155_o = flagssr[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:47  */
  assign n1156_o = $unsigned(n1155_o) < $unsigned(ipl_nr);
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:64  */
  assign n1158_o = ipl_nr == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:55  */
  assign n1159_o = n1156_o | n1158_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:72  */
  assign n1160_o = n1159_o | make_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:90  */
  assign n1161_o = n1160_o | make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1043:35  */
  assign n1162_o = ~stop;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1043:25  */
  assign n1165_o = n1162_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:25  */
  assign n1167_o = n1161_o ? 1'b0 : n1165_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1041:25  */
  assign n1170_o = n1161_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:17  */
  assign n1172_o = n1154_o ? n1167_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:17  */
  assign n1176_o = n1154_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1039:17  */
  assign n1179_o = n1154_o ? n1170_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:28  */
  assign n1182_o = setstate == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:54  */
  assign n1184_o = next_micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:34  */
  assign n1185_o = n1182_o & n1184_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:79  */
  assign n1186_o = ~set_direct_data;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:60  */
  assign n1187_o = n1185_o & n1186_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:104  */
  assign n1188_o = ~exec_write_back;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:118  */
  assign n1190_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:137  */
  assign n1191_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:124  */
  assign n1192_o = n1190_o & n1191_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:109  */
  assign n1193_o = n1188_o | n1192_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:84  */
  assign n1194_o = n1187_o & n1193_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1048:17  */
  assign n1197_o = n1194_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1052:27  */
  assign n1199_o = ~ipl;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1082:59  */
  assign n1201_o = memmask[3:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1082:71  */
  assign n1203_o = {n1201_o, 2'b11};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1083:59  */
  assign n1204_o = memread[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1083:82  */
  assign n1205_o = memmaskmux[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1083:71  */
  assign n1206_o = {n1204_o, n1205_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1087:48  */
  assign n1207_o = exec[57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1089:51  */
  assign n1208_o = exec[63];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1091:54  */
  assign n1210_o = state == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1091:60  */
  assign n1211_o = n1210_o | tg68_pc_brw;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1091:90  */
  assign n1212_o = ~stop;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1091:82  */
  assign n1213_o = n1211_o & n1212_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1091:41  */
  assign n1214_o = n1213_o ? tg68_pc_add : tg68_pc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1089:41  */
  assign n1215_o = n1208_o ? addr : n1214_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1087:41  */
  assign n1216_o = n1207_o ? data_read : n1215_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1081:33  */
  assign n1217_o = clkena_in ? n1216_o : tg68_pc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1081:33  */
  assign n1218_o = clkena_in ? n1203_o : memmask;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1081:33  */
  assign n1219_o = clkena_in ? n1206_o : memread;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1109:53  */
  assign n1220_o = ~trap_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1110:68  */
  assign n1221_o = berr | make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1109:41  */
  assign n1223_o = n1220_o ? n1221_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1115:71  */
  assign n1224_o = ~setinterrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1115:67  */
  assign n1225_o = stop & n1224_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1115:58  */
  assign n1226_o = set_stop | n1225_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1128:75  */
  assign n1228_o = {5'b00011, ipl_nr};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1124:49  */
  assign n1231_o = make_berr ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1124:49  */
  assign n1234_o = make_berr ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1124:49  */
  assign n1235_o = make_berr ? ripl_nr : ipl_nr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1124:49  */
  assign n1236_o = make_berr ? ipl_vec : n1228_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1122:49  */
  assign n1238_o = make_trace ? 1'b0 : n1231_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1122:49  */
  assign n1242_o = make_trace ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1122:49  */
  assign n1245_o = make_trace ? 1'b0 : n1234_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1122:49  */
  assign n1247_o = make_trace ? ripl_nr : n1235_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1122:49  */
  assign n1248_o = make_trace ? ipl_vec : n1236_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1116:41  */
  assign n1249_o = setinterrupt ? n1238_o : trap_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1116:41  */
  assign n1250_o = setinterrupt ? n1242_o : trap_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1116:41  */
  assign n1251_o = setinterrupt ? n1245_o : trap_interrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1116:41  */
  assign n1253_o = setinterrupt ? 1'b0 : n1223_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1254_o = n1457_o ? n1247_o : ripl_nr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1116:41  */
  assign n1255_o = setinterrupt ? n1248_o : ipl_vec;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1132:55  */
  assign n1257_o = micro_state == 7'b0110011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1132:80  */
  assign n1258_o = ~ipl_autovector;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1132:62  */
  assign n1259_o = n1257_o & n1258_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1133:74  */
  assign n1260_o = last_data_read[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1132:41  */
  assign n1261_o = n1259_o ? n1260_o : n1255_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1135:49  */
  assign n1263_o = state == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1136:75  */
  assign n1264_o = data_read[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1265_o = n1439_o ? tg68_pc : last_opc_pc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1266_o = n1440_o ? n1264_o : last_opc_read;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1144:53  */
  assign n1267_o = opcode[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1144:65  */
  assign n1269_o = n1267_o == 8'b00000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1144:86  */
  assign n1270_o = opcode[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1144:98  */
  assign n1272_o = n1270_o == 8'b11111111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1144:77  */
  assign n1273_o = n1269_o | n1272_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1144:110  */
  assign n1274_o = n1273_o | data_is_source;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1144:41  */
  assign n1276_o = n1274_o ? 1'b1 : tg68_pc_word;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1139:41  */
  assign n1278_o = setopcode ? 1'b0 : n1276_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1139:41  */
  assign n1280_o = setopcode ? 1'b0 : n1249_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1139:41  */
  assign n1282_o = setopcode ? 1'b0 : n1250_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1139:41  */
  assign n1284_o = setopcode ? 1'b0 : n1251_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1148:48  */
  assign n1285_o = exec[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1152:84  */
  assign n1286_o = {26'b0, bf_width};  //  uext
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1152:84  */
  assign n1287_o = bf_full_offset + n1286_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1152:93  */
  assign n1289_o = n1287_o + 32'b00000000000000000000000000000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1290_o = n1466_o ? bf_width : alu_width;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1291_o = n1467_o ? bf_shift : alu_bf_shift;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1292_o = n1468_o ? n1289_o : alu_bf_ffo_offset;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1293_o = n1469_o ? bf_loffset : alu_bf_loffset;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1155:62  */
  assign n1294_o = setstate[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1155:50  */
  assign n1295_o = ~n1294_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1155:93  */
  assign n1296_o = setstate[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1155:81  */
  assign n1297_o = ~n1296_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1155:77  */
  assign n1298_o = pcbase & n1297_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1155:66  */
  assign n1299_o = n1295_o | n1298_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1156:58  */
  assign n1300_o = setstate[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1156:67  */
  assign n1301_o = ~pcbase;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1156:89  */
  assign n1302_o = setstate[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1156:78  */
  assign n1303_o = n1301_o | n1302_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1156:62  */
  assign n1304_o = n1300_o & n1303_o;
  assign n1306_o = {n1299_o, n1304_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1157:41  */
  assign n1307_o = interrupt ? 2'b11 : n1306_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1161:49  */
  assign n1309_o = state == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1163:55  */
  assign n1311_o = setstate == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1163:77  */
  assign n1312_o = ~setaddrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1163:61  */
  assign n1313_o = n1311_o & n1312_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1163:82  */
  assign n1314_o = n1313_o & write_back;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1163:41  */
  assign n1316_o = n1314_o ? 1'b1 : exec_write_back;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1161:41  */
  assign n1318_o = n1309_o ? 1'b0 : n1316_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:50  */
  assign n1320_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:69  */
  assign n1321_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:56  */
  assign n1322_o = n1320_o & n1321_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:74  */
  assign n1323_o = n1322_o & write_back;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:105  */
  assign n1325_o = setstate != 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:93  */
  assign n1326_o = n1323_o & n1325_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:127  */
  assign n1328_o = set_rot_cnt != 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:113  */
  assign n1329_o = n1326_o | n1328_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:164  */
  assign n1330_o = ~interrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:151  */
  assign n1331_o = stop & n1330_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:138  */
  assign n1332_o = n1329_o | n1331_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:181  */
  assign n1333_o = set_exec[31];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:170  */
  assign n1334_o = n1332_o | n1333_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1170:59  */
  assign n1335_o = execopc & exec_write_back;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1178:60  */
  assign n1338_o = setstate == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1181:59  */
  assign n1339_o = exec[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1185:58  */
  assign n1340_o = set[73];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1190:67  */
  assign n1342_o = set_datatype == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1190:85  */
  assign n1343_o = setstate[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1190:73  */
  assign n1344_o = n1342_o & n1343_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1193:63  */
  assign n1345_o = set[72];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1193:57  */
  assign n1348_o = n1345_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1190:49  */
  assign n1351_o = n1344_o ? 6'b101111 : 6'b100111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1190:49  */
  assign n1354_o = n1344_o ? 6'b101111 : 6'b100111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1190:49  */
  assign n1356_o = n1344_o ? n1348_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1185:49  */
  assign n1358_o = n1340_o ? 6'b100001 : n1351_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1185:49  */
  assign n1360_o = n1340_o ? 6'b100001 : n1354_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1185:49  */
  assign n1362_o = n1340_o ? 1'b0 : n1356_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1181:49  */
  assign n1363_o = n1339_o ? set_memmask : n1358_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1181:49  */
  assign n1364_o = n1339_o ? set_memmask : n1360_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1181:49  */
  assign n1365_o = n1339_o ? set_oddout : n1362_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1178:49  */
  assign n1367_o = n1338_o ? 6'b111111 : n1363_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1178:49  */
  assign n1369_o = n1338_o ? 6'b111111 : n1364_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1178:49  */
  assign n1370_o = n1338_o ? oddout : n1365_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1170:41  */
  assign n1371_o = n1335_o ? 2'b01 : n1307_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1170:41  */
  assign n1373_o = n1335_o ? 2'b11 : setstate;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1170:41  */
  assign n1375_o = n1335_o ? 1'b0 : setaddrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1170:41  */
  assign n1376_o = n1335_o ? wbmemmask : n1367_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1170:41  */
  assign n1377_o = n1335_o ? wbmemmask : n1369_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1170:41  */
  assign n1378_o = n1335_o ? oddout : n1370_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:41  */
  assign n1379_o = n1334_o ? n1307_o : n1371_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:41  */
  assign n1381_o = n1334_o ? 2'b01 : n1373_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:41  */
  assign n1383_o = n1334_o ? 1'b0 : n1375_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:41  */
  assign n1385_o = n1334_o ? 6'b111111 : n1376_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:41  */
  assign n1386_o = n1334_o ? wbmemmask : n1377_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1166:41  */
  assign n1387_o = n1334_o ? oddout : n1378_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1209:78  */
  assign n1388_o = set_writepcbig | writepcbig;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1205:41  */
  assign n1390_o = decodeopc ? 1'b0 : n1388_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1391_o = n1449_o ? set_rot_bits : rot_bits;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1211:65  */
  assign n1392_o = exec[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1211:58  */
  assign n1393_o = decodeopc | n1392_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1211:92  */
  assign n1395_o = rot_cnt != 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1211:82  */
  assign n1396_o = n1393_o | n1395_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1397_o = n1450_o ? set_rot_cnt : rot_cnt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1217:55  */
  assign n1398_o = setstate[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1217:86  */
  assign n1399_o = set[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1217:79  */
  assign n1400_o = ea_only & n1399_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1217:63  */
  assign n1401_o = n1398_o | n1400_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1217:41  */
  assign n1403_o = n1401_o ? 1'b0 : suppress_base;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1215:41  */
  assign n1405_o = set_suppress_base ? 1'b1 : n1403_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1221:57  */
  assign n1406_o = state[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1224:75  */
  assign n1407_o = data_read[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1221:49  */
  assign n1408_o = n1406_o ? last_opc_read : n1407_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1409_o = n1443_o ? n1408_o : brief;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1228:66  */
  assign n1410_o = ~berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1228:58  */
  assign n1411_o = setopcode & n1410_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1229:57  */
  assign n1413_o = state == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1230:76  */
  assign n1414_o = data_read[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1229:49  */
  assign n1415_o = n1413_o ? n1414_o : last_opc_read;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1229:49  */
  assign n1416_o = n1413_o ? tg68_pc : last_opc_pc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1237:64  */
  assign n1417_o = setinterrupt | setopcode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1242:68  */
  assign n1418_o = setnextpass | regdirectsource;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1242:49  */
  assign n1420_o = n1418_o ? 1'b1 : nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1237:41  */
  assign n1422_o = n1417_o ? 16'b0100111001110001 : opcode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1237:41  */
  assign n1424_o = n1417_o ? 1'b0 : n1420_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1228:41  */
  assign n1425_o = n1411_o ? n1415_o : n1422_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1426_o = n1438_o ? n1416_o : exe_pc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1228:41  */
  assign n1428_o = n1411_o ? 1'b0 : n1424_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1247:58  */
  assign n1429_o = decodeopc | interrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1430_o = n1454_o ? flagssr : trap_sr;
  assign n1431_o = n9523_o[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1432_o = clkena_lw ? n1379_o : n1431_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1433_o = clkena_lw ? n1381_o : state;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1434_o = clkena_lw ? set_datatype : exe_datatype;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1435_o = clkena_lw ? n1383_o : addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1436_o = clkena_lw ? n1425_o : opcode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1437_o = clkena_lw ? opcode : exe_opcode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1438_o = clkena_lw & n1411_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1439_o = clkena_lw & n1263_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1440_o = clkena_lw & n1263_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1441_o = clkena_lw ? n1428_o : nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1442_o = clkena_lw ? n1278_o : tg68_pc_word;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1443_o = clkena_lw & getbrief;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1444_o = clkena_lw ? n1318_o : exec_write_back;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1445_o = clkena_lw ? n1390_o : writepcbig;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1446_o = clkena_lw ? setopcode : decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1447_o = clkena_lw ? setexecopc : execopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1448_o = clkena_lw ? setendopc : endopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1449_o = clkena_lw & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1450_o = clkena_lw & n1396_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1451_o = clkena_lw ? n1280_o : trap_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1452_o = clkena_lw ? n1282_o : trap_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1453_o = clkena_lw ? n1284_o : trap_interrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1454_o = clkena_lw & n1429_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1455_o = clkena_lw ? n1253_o : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1456_o = clkena_lw ? n1226_o : stop;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1457_o = clkena_lw & setinterrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1458_o = clkena_lw ? n1261_o : ipl_vec;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1459_o = clkena_lw ? setinterrupt : interrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1460_o = clkena_lw ? n1405_o : suppress_base;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1461_o = clkena_lw ? n1385_o : n1218_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1463_o = clkena_lw ? 4'b1111 : n1219_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1464_o = clkena_lw ? n1386_o : wbmemmask;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1465_o = clkena_lw ? n1387_o : oddout;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1466_o = clkena_lw & n1285_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1467_o = clkena_lw & n1285_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1468_o = clkena_lw & n1285_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1095:33  */
  assign n1469_o = clkena_lw & n1285_o;
  assign n1470_o = n9523_o[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1471_o = reset ? n1470_o : n1432_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1473_o = reset ? 32'b00000000000000000000000000000100 : n1217_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1475_o = reset ? 2'b01 : n1433_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1476_o = reset ? exe_datatype : n1434_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1478_o = reset ? 1'b0 : n1435_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1480_o = reset ? 16'b0010111001111001 : n1436_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1481_o = reset ? exe_opcode : n1437_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1482_o = reset ? exe_pc : n1426_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1483_o = reset ? last_opc_pc : n1265_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1485_o = reset ? 16'b0100111011111001 : n1266_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1486_o = reset ? nextpass : n1441_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1488_o = reset ? 1'b0 : n1442_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1489_o = reset ? brief : n1409_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1491_o = reset ? 1'b0 : n1444_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1493_o = reset ? 1'b0 : n1445_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1495_o = reset ? 1'b0 : n1446_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1497_o = reset ? 1'b0 : n1447_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1499_o = reset ? 1'b0 : n1448_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1500_o = reset ? rot_bits : n1391_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1502_o = reset ? 6'b000001 : n1397_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1504_o = reset ? 1'b0 : n1451_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1506_o = reset ? 1'b0 : n1452_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1508_o = reset ? 1'b0 : n1453_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1509_o = reset ? trap_sr : n1430_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1511_o = reset ? 1'b0 : n1455_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1513_o = reset ? 1'b0 : n1456_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1514_o = reset ? ripl_nr : n1254_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1515_o = reset ? ipl_vec : n1458_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1517_o = reset ? 1'b0 : n1459_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1519_o = reset ? 1'b0 : n1460_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1521_o = reset ? 6'b111111 : n1461_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1522_o = reset ? memread : n1463_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1523_o = reset ? wbmemmask : n1464_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1524_o = reset ? oddout : n1465_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1525_o = reset ? alu_width : n1290_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1526_o = reset ? alu_bf_shift : n1291_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1527_o = reset ? alu_bf_ffo_offset : n1292_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1054:25  */
  assign n1528_o = reset ? alu_bf_loffset : n1293_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1258:54  */
  assign n1569_o = set_pcbase | pcbase;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1259:60  */
  assign n1570_o = state[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1259:81  */
  assign n1571_o = ~movem_run;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1259:68  */
  assign n1572_o = n1570_o & n1571_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1259:51  */
  assign n1573_o = setexecopc | n1572_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1259:33  */
  assign n1575_o = n1573_o ? 1'b0 : n1569_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1257:25  */
  assign n1576_o = clkena_lw ? n1575_o : pcbase;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1255:25  */
  assign n1578_o = reset ? 1'b1 : n1576_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1265:54  */
  assign n1579_o = set[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1265:70  */
  assign n1580_o = set[85];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1265:64  */
  assign n1581_o = n1579_o | n1580_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1266:58  */
  assign n1584_o = set[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1266:73  */
  assign n1585_o = set[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1266:67  */
  assign n1586_o = n1584_o | n1585_o;
  assign n1587_o = set[88:87];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1268:52  */
  assign n1588_o = set[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1268:67  */
  assign n1589_o = set[48];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1268:61  */
  assign n1590_o = n1588_o | n1589_o;
  assign n1591_o = set[84:49];
  assign n1592_o = set[47:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1270:58  */
  assign n1593_o = set_exec | set;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1271:67  */
  assign n1594_o = set_exec[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1271:83  */
  assign n1595_o = set[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1271:77  */
  assign n1596_o = n1594_o | n1595_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1271:99  */
  assign n1597_o = set[85];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1271:93  */
  assign n1598_o = n1596_o | n1597_o;
  assign n1600_o = n1593_o[84:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1272:71  */
  assign n1601_o = set_exec[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1272:86  */
  assign n1602_o = set[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1272:80  */
  assign n1603_o = n1601_o | n1602_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1272:101  */
  assign n1604_o = set[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1272:95  */
  assign n1605_o = n1603_o | n1604_o;
  assign n1606_o = n1593_o[88:87];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1269:33  */
  assign n1608_o = setexecopc ? set_exec_tas : 1'b0;
  assign n1610_o = {n1606_o, n1605_o, n1598_o, n1600_o};
  assign n1611_o = {n1587_o, n1586_o, n1581_o, n1591_o, n1590_o, n1592_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1275:56  */
  assign n1613_o = set[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1275:69  */
  assign n1614_o = n1613_o | setopcode;
  assign n1615_o = n1610_o[88:72];
  assign n1616_o = n1611_o[88:72];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1269:33  */
  assign n1617_o = setexecopc ? n1615_o : n1616_o;
  assign n1618_o = n1610_o[70:0];
  assign n1619_o = n1611_o[70:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1269:33  */
  assign n1620_o = setexecopc ? n1618_o : n1619_o;
  assign n1622_o = {n1617_o, n1614_o, n1620_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1285:26  */
  assign n1630_o = sndopc[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1286:48  */
  assign n1631_o = reg_qa[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1286:41  */
  assign n1633_o = {1'b0, n1631_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1288:48  */
  assign n1634_o = sndopc[10:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1288:41  */
  assign n1636_o = {1'b0, n1634_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1290:26  */
  assign n1638_o = sndopc[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1294:61  */
  assign n1639_o = sndopc[10:6];
  assign n1641_o = n1640_o[31:5];
  assign n1642_o = {n1641_o, n1639_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1290:17  */
  assign n1643_o = n1638_o ? reg_qa : n1642_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1298:26  */
  assign n1645_o = sndopc[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1299:55  */
  assign n1646_o = reg_qb[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1299:67  */
  assign n1648_o = n1646_o - 5'b00001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1301:55  */
  assign n1649_o = sndopc[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1301:67  */
  assign n1651_o = n1649_o - 5'b00001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1298:17  */
  assign n1652_o = n1645_o ? n1648_o : n1651_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1303:37  */
  assign n1653_o = bf_width + bf_offset;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1304:43  */
  assign n1654_o = bf_bhits[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1304:31  */
  assign n1655_o = ~n1654_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1308:26  */
  assign n1656_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1308:39  */
  assign n1658_o = n1656_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1309:41  */
  assign n1660_o = 6'b100000 - bf_shift;
  assign n1663_o = n1660_o[4:0];
  assign n1664_o = bf_shift[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1308:17  */
  assign n1665_o = n1658_o ? n1663_o : n1664_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1315:26  */
  assign n1666_o = opcode[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1315:38  */
  assign n1668_o = n1666_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1316:34  */
  assign n1669_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1316:47  */
  assign n1671_o = n1669_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1317:53  */
  assign n1673_o = bf_bhits + 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1319:47  */
  assign n1675_o = 6'b011111 - bf_bhits;
  assign n1678_o = n1673_o[4:0];
  assign n1679_o = n1675_o[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1316:25  */
  assign n1680_o = n1671_o ? n1678_o : n1679_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1323:34  */
  assign n1681_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1323:47  */
  assign n1683_o = n1681_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1324:69  */
  assign n1684_o = bf_bhits[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1324:60  */
  assign n1686_o = {3'b000, n1684_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1324:53  */
  assign n1688_o = 6'b011001 + n1686_o;
  assign n1690_o = n1688_o[4:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1327:66  */
  assign n1691_o = bf_bhits[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1327:57  */
  assign n1693_o = 3'b111 - n1691_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1327:50  */
  assign n1695_o = {3'b000, n1693_o};
  assign n1696_o = {1'b0, n1690_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1323:25  */
  assign n1697_o = n1683_o ? n1696_o : n1695_o;
  assign n1699_o = n1633_o[4:3];
  assign n1700_o = n1636_o[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1285:17  */
  assign n1701_o = n1630_o ? n1699_o : n1700_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1315:17  */
  assign n1702_o = n1668_o ? n1701_o : 2'b00;
  assign n1703_o = n1633_o[5];
  assign n1704_o = n1636_o[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1285:17  */
  assign n1705_o = n1630_o ? n1703_o : n1704_o;
  assign n1706_o = n1633_o[2:0];
  assign n1707_o = n1636_o[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1285:17  */
  assign n1708_o = n1630_o ? n1706_o : n1707_o;
  assign n1709_o = {1'b0, n1680_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1315:17  */
  assign n1710_o = n1668_o ? n1709_o : n1697_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1332:30  */
  assign n1711_o = bf_bhits[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1333:25  */
  assign n1713_o = n1711_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1335:25  */
  assign n1715_o = n1711_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1337:25  */
  assign n1717_o = n1711_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1339:25  */
  assign n1719_o = n1711_o == 3'b011;
  assign n1720_o = {n1719_o, n1717_o, n1715_o, n1713_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1332:17  */
  always @*
    case (n1720_o)
      4'b1000: n1726_o = 6'b100001;
      4'b0100: n1726_o = 6'b100011;
      4'b0010: n1726_o = 6'b100111;
      4'b0001: n1726_o = 6'b101111;
      default: n1726_o = 6'b100000;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1344:28  */
  assign n1728_o = setstate == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1344:17  */
  assign n1730_o = n1728_o ? 6'b100111 : n1726_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1354:24  */
  assign n1734_o = exec[17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1355:59  */
  assign n1735_o = last_data_read[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1355:41  */
  assign n1736_o = flagssr & n1735_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1356:27  */
  assign n1737_o = exec[18];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1357:59  */
  assign n1738_o = last_data_read[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1357:41  */
  assign n1739_o = flagssr ^ n1738_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1358:27  */
  assign n1740_o = exec[19];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1359:58  */
  assign n1741_o = last_data_read[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1359:41  */
  assign n1742_o = flagssr | n1741_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1361:39  */
  assign n1743_o = op2out[15:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1358:17  */
  assign n1744_o = n1740_o ? n1742_o : n1743_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1356:17  */
  assign n1745_o = n1737_o ? n1739_o : n1744_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1354:17  */
  assign n1746_o = n1734_o ? n1736_o : n1745_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1373:62  */
  assign n1749_o = flagssr[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1374:47  */
  assign n1750_o = set[41];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1375:59  */
  assign n1751_o = ~svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1374:41  */
  assign n1752_o = n1750_o ? n1751_o : presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1372:33  */
  assign n1753_o = setopcode ? n1749_o : make_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1371:25  */
  assign n1754_o = n1841_o ? n1752_o : svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1380:50  */
  assign n1755_o = trap_berr | trap_illegal;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1380:70  */
  assign n1756_o = n1755_o | trap_addr_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1380:93  */
  assign n1757_o = n1756_o | trap_priv;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1380:110  */
  assign n1758_o = n1757_o | trap_1010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1380:127  */
  assign n1759_o = n1758_o | trap_1111;
  assign n1761_o = flagssr[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1380:33  */
  assign n1762_o = n1759_o ? 1'b0 : n1761_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1380:33  */
  assign n1764_o = n1759_o ? 1'b0 : n1753_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1384:39  */
  assign n1765_o = set[41];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1385:54  */
  assign n1766_o = ~presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1386:55  */
  assign n1767_o = ~presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1387:50  */
  assign n1768_o = ~presvmode;
  assign n1769_o = n9523_o[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1384:33  */
  assign n1770_o = n1765_o ? n1768_o : n1769_o;
  assign n1771_o = flagssr[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1384:33  */
  assign n1772_o = n1765_o ? n1767_o : n1771_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1371:25  */
  assign n1773_o = n1842_o ? n1766_o : presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1389:47  */
  assign n1775_o = micro_state == 7'b0110110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1389:33  */
  assign n1777_o = n1775_o ? 1'b0 : n1762_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1392:60  */
  assign n1779_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1392:51  */
  assign n1780_o = trap_trace & n1779_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1392:33  */
  assign n1782_o = n1780_o ? 1'b0 : n1764_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1395:40  */
  assign n1783_o = exec[59];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1395:55  */
  assign n1784_o = n1783_o | set_stop;
  assign n1786_o = flagssr[4:0];
  assign n1787_o = flagssr[6];
  assign n1788_o = {n1777_o, n1787_o, n1772_o, n1786_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1398:50  */
  assign n1790_o = interrupt & trap_interrupt;
  assign n1791_o = data_read[10:8];
  assign n1792_o = n1788_o[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1395:33  */
  assign n1793_o = n1784_o ? n1791_o : n1792_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1398:33  */
  assign n1794_o = n1790_o ? ripl_nr : n1793_o;
  assign n1795_o = data_read[15:11];
  assign n1796_o = n1788_o[7:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1395:33  */
  assign n1797_o = n1784_o ? n1795_o : n1796_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1401:40  */
  assign n1798_o = exec[52];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1403:54  */
  assign n1799_o = srin[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1404:43  */
  assign n1800_o = exec[35];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1405:57  */
  assign n1801_o = flagssr[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1404:33  */
  assign n1802_o = n1800_o ? n1801_o : n1770_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1401:33  */
  assign n1803_o = n1798_o ? n1799_o : n1802_o;
  assign n1804_o = {n1797_o, n1794_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1407:33  */
  assign n1807_o = interrupt ? 1'b1 : n1803_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1410:39  */
  assign n1808_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1410:42  */
  assign n1809_o = ~n1808_o;
  assign n1812_o = srin[4];
  assign n1813_o = n1804_o[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1401:33  */
  assign n1814_o = n1798_o ? n1812_o : n1813_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1410:33  */
  assign n1815_o = n1809_o ? 1'b0 : n1814_o;
  assign n1816_o = srin[6];
  assign n1817_o = n1804_o[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1401:33  */
  assign n1818_o = n1798_o ? n1816_o : n1817_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1410:33  */
  assign n1819_o = n1809_o ? 1'b0 : n1818_o;
  assign n1826_o = srin[7];
  assign n1827_o = n1804_o[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1401:33  */
  assign n1828_o = n1798_o ? n1826_o : n1827_o;
  assign n1829_o = srin[5];
  assign n1830_o = n1804_o[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1401:33  */
  assign n1831_o = n1798_o ? n1829_o : n1830_o;
  assign n1833_o = srin[2:0];
  assign n1834_o = n1804_o[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1401:33  */
  assign n1835_o = n1798_o ? n1833_o : n1834_o;
  assign n1836_o = n9523_o[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1371:25  */
  assign n1837_o = clkena_lw ? n1807_o : n1836_o;
  assign n1838_o = {n1828_o, n1819_o, n1831_o, n1815_o, 1'b0, n1835_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1371:25  */
  assign n1839_o = clkena_lw ? n1838_o : flagssr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1371:25  */
  assign n1840_o = clkena_lw ? n1782_o : make_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1371:25  */
  assign n1841_o = clkena_lw & setopcode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1371:25  */
  assign n1842_o = clkena_lw & n1765_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1365:25  */
  assign n1843_o = reset ? 1'b1 : n1837_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1365:25  */
  assign n1845_o = reset ? 8'b00100111 : n1839_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1365:25  */
  assign n1847_o = reset ? 1'b0 : n1840_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1365:25  */
  assign n1849_o = reset ? 1'b1 : n1754_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1365:25  */
  assign n1851_o = reset ? 1'b1 : n1773_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1447:39  */
  assign n1861_o = opcode[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1489:27  */
  assign n1863_o = rot_cnt != 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1490:47  */
  assign n1865_o = rot_cnt - 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1489:17  */
  assign n1867_o = n1863_o ? n1865_o : 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1501:28  */
  assign n1873_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1502:25  */
  assign n1875_o = n1873_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1503:25  */
  assign n1877_o = n1873_o == 2'b01;
  assign n1878_o = {n1877_o, n1875_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1501:17  */
  always @*
    case (n1878_o)
      2'b10: n1882_o = 2'b01;
      2'b01: n1882_o = 2'b00;
      default: n1882_o = 2'b10;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1507:32  */
  assign n1883_o = execopc & exec_write_back;
  assign n1885_o = n1870_o[83];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1507:17  */
  assign n1886_o = n1883_o ? 1'b1 : n1885_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1511:34  */
  assign n1889_o = interrupt & trap_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1513:37  */
  assign n1890_o = ~presvmode;
  assign n1892_o = n1870_o[41];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1511:17  */
  assign n1893_o = n1899_o ? 1'b1 : n1892_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1511:17  */
  assign n1896_o = n1889_o ? 2'b01 : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1511:17  */
  assign n1899_o = n1889_o & n1890_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1511:17  */
  assign n1904_o = n1889_o ? 7'b0110011 : 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:42  */
  assign n1906_o = ~trapd;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:33  */
  assign n1907_o = trapmake & n1906_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1519:31  */
  assign n1908_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1519:59  */
  assign n1909_o = trap_trapv | set_z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1519:85  */
  assign n1910_o = exec[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1519:78  */
  assign n1911_o = n1909_o | n1910_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1519:39  */
  assign n1912_o = n1908_o & n1911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1519:25  */
  assign n1915_o = n1912_o ? 7'b0110010 : 7'b0110011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1524:46  */
  assign n1916_o = ~use_vbr_stackframe;
  assign n1918_o = n1870_o[25];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:17  */
  assign n1919_o = n1926_o ? 1'b1 : n1918_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1528:37  */
  assign n1920_o = ~presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:17  */
  assign n1922_o = n1927_o ? 1'b1 : n1893_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:17  */
  assign n1924_o = n1907_o ? 2'b01 : n1896_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:17  */
  assign n1926_o = n1907_o & n1916_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:17  */
  assign n1927_o = n1907_o & n1920_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1518:17  */
  assign n1930_o = n1907_o ? n1915_o : n1904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1533:31  */
  assign n1932_o = micro_state == 7'b0100111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1533:55  */
  assign n1933_o = interrupt & trap_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1533:37  */
  assign n1934_o = n1932_o | n1933_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1535:50  */
  assign n1935_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1535:43  */
  assign n1936_o = trap_trace & n1935_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1535:25  */
  assign n1939_o = n1936_o ? 7'b0110010 : 7'b0110011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1545:37  */
  assign n1940_o = ~presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1533:17  */
  assign n1942_o = n1945_o ? 1'b1 : n1922_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1533:17  */
  assign n1944_o = n1934_o ? 2'b01 : n1924_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1533:17  */
  assign n1945_o = n1934_o & n1940_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1533:17  */
  assign n1946_o = n1934_o ? n1939_o : n1930_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1550:24  */
  assign n1948_o = micro_state == 7'b0100111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1550:51  */
  assign n1949_o = interrupt & trap_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1550:31  */
  assign n1950_o = n1948_o | n1949_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1551:24  */
  assign n1951_o = ~presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1550:9  */
  assign n1953_o = n1956_o ? 1'b1 : n1942_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1550:9  */
  assign n1955_o = n1950_o ? 2'b01 : n1944_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1550:9  */
  assign n1956_o = n1950_o & n1951_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1557:46  */
  assign n1957_o = flagssr[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1557:49  */
  assign n1958_o = n1957_o != presvmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1557:35  */
  assign n1959_o = setexecopc & n1958_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1557:17  */
  assign n1961_o = n1959_o ? 1'b1 : n1953_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1563:34  */
  assign n1962_o = interrupt & trap_interrupt;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1563:17  */
  assign n1965_o = n1962_o ? 2'b10 : n1955_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1563:17  */
  assign n1966_o = n1962_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1563:17  */
  assign n1968_o = n1962_o ? 7'b0100111 : n1946_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:23  */
  assign n1969_o = set[41];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:17  */
  assign n1974_o = n1969_o ? 1'b1 : 1'b0;
  assign n1976_o = {1'b1, 1'b1};
  assign n1977_o = n1870_o[66:65];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:17  */
  assign n1978_o = n1969_o ? n1976_o : n1977_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1576:27  */
  assign n1981_o = ~ea_only;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1576:39  */
  assign n1982_o = set[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1576:32  */
  assign n1983_o = n1981_o & n1982_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1576:17  */
  assign n1985_o = n1983_o ? 2'b10 : n1965_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1582:28  */
  assign n1986_o = setstate[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1582:52  */
  assign n1987_o = set_datatype[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1582:36  */
  assign n1988_o = n1986_o & n1987_o;
  assign n1990_o = n1870_o[73];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1582:17  */
  assign n1991_o = n1988_o ? 1'b1 : n1990_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:38  */
  assign n1994_o = ea_build_now & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:64  */
  assign n1995_o = exec[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:57  */
  assign n1996_o = n1994_o | n1995_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:36  */
  assign n1997_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1591:50  */
  assign n1999_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1593:58  */
  assign n2001_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1593:70  */
  assign n2003_o = n2001_o == 3'b111;
  assign n2005_o = n1870_o[50];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1591:41  */
  assign n2006_o = n2010_o ? 1'b1 : n2005_o;
  assign n2007_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1591:41  */
  assign n2008_o = n1999_o ? 1'b1 : n2007_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1591:41  */
  assign n2010_o = n1999_o & n2003_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1597:50  */
  assign n2011_o = opcode[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1599:58  */
  assign n2013_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1599:70  */
  assign n2015_o = n2013_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1597:41  */
  assign n2017_o = n2020_o ? 1'b1 : n2006_o;
  assign n2018_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1597:41  */
  assign n2019_o = n2011_o ? 1'b1 : n2018_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1597:41  */
  assign n2020_o = n2011_o & n2015_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1588:33  */
  assign n2022_o = n1997_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1588:43  */
  assign n2024_o = n1997_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1588:43  */
  assign n2025_o = n2022_o | n2024_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1588:49  */
  assign n2027_o = n1997_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1588:49  */
  assign n2028_o = n2025_o | n2027_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1603:33  */
  assign n2030_o = n1997_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1605:33  */
  assign n2032_o = n1997_o == 3'b110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:52  */
  assign n2033_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1610:49  */
  assign n2035_o = n2033_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1612:49  */
  assign n2038_o = n2033_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1615:49  */
  assign n2041_o = n2033_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1620:49  */
  assign n2044_o = n2033_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1629:68  */
  assign n2046_o = datatype == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1629:57  */
  assign n2048_o = n2046_o ? 1'b1 : n1991_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1626:49  */
  assign n2050_o = n2033_o == 3'b100;
  assign n2051_o = {n2050_o, n2044_o, n2041_o, n2038_o, n2035_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2054_o = 1'b1;
      5'b01000: n2054_o = 1'b0;
      5'b00100: n2054_o = 1'b0;
      5'b00010: n2054_o = 1'b0;
      5'b00001: n2054_o = 1'b0;
      default: n2054_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2057_o = 1'b0;
      5'b01000: n2057_o = 1'b1;
      5'b00100: n2057_o = 1'b0;
      5'b00010: n2057_o = 1'b0;
      5'b00001: n2057_o = 1'b0;
      default: n2057_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2060_o = 1'b1;
      5'b01000: n2060_o = 1'b0;
      5'b00100: n2060_o = 1'b0;
      5'b00010: n2060_o = 1'b0;
      5'b00001: n2060_o = 1'b0;
      default: n2060_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2064_o = 1'b0;
      5'b01000: n2064_o = 1'b1;
      5'b00100: n2064_o = 1'b1;
      5'b00010: n2064_o = 1'b0;
      5'b00001: n2064_o = 1'b0;
      default: n2064_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2068_o = 1'b0;
      5'b01000: n2068_o = 1'b1;
      5'b00100: n2068_o = 1'b1;
      5'b00010: n2068_o = 1'b0;
      5'b00001: n2068_o = 1'b0;
      default: n2068_o = 1'b0;
    endcase
  assign n2069_o = n1870_o[22];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2070_o = n2069_o;
      5'b01000: n2070_o = 1'b1;
      5'b00100: n2070_o = 1'b1;
      5'b00010: n2070_o = n2069_o;
      5'b00001: n2070_o = n2069_o;
      default: n2070_o = n2069_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2071_o = n2048_o;
      5'b01000: n2071_o = n1991_o;
      5'b00100: n2071_o = n1991_o;
      5'b00010: n2071_o = 1'b1;
      5'b00001: n2071_o = n1991_o;
      default: n2071_o = n1991_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1609:41  */
  always @*
    case (n2051_o)
      5'b10000: n2076_o = n1968_o;
      5'b01000: n2076_o = 7'b0000101;
      5'b00100: n2076_o = 7'b0000100;
      5'b00010: n2076_o = 7'b0000010;
      5'b00001: n2076_o = 7'b0000010;
      default: n2076_o = n1968_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1608:33  */
  assign n2078_o = n1997_o == 3'b111;
  assign n2079_o = {n2078_o, n2032_o, n2030_o, n2028_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2082_o = n2054_o;
      4'b0100: n2082_o = 1'b0;
      4'b0010: n2082_o = 1'b0;
      4'b0001: n2082_o = 1'b1;
      default: n2082_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2085_o = n2057_o;
      4'b0100: n2085_o = 1'b1;
      4'b0010: n2085_o = 1'b0;
      4'b0001: n2085_o = 1'b0;
      default: n2085_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2087_o = n2060_o;
      4'b0100: n2087_o = 1'b0;
      4'b0010: n2087_o = 1'b0;
      4'b0001: n2087_o = 1'b0;
      default: n2087_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2089_o = n2064_o;
      4'b0100: n2089_o = 1'b0;
      4'b0010: n2089_o = 1'b0;
      4'b0001: n2089_o = 1'b0;
      default: n2089_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2091_o = n2068_o;
      4'b0100: n2091_o = 1'b0;
      4'b0010: n2091_o = 1'b0;
      4'b0001: n2091_o = 1'b0;
      default: n2091_o = 1'b0;
    endcase
  assign n2092_o = n1870_o[22];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2093_o = n2070_o;
      4'b0100: n2093_o = n2092_o;
      4'b0010: n2093_o = n2092_o;
      4'b0001: n2093_o = n2092_o;
      default: n2093_o = n2092_o;
    endcase
  assign n2094_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2095_o = n2094_o;
      4'b0100: n2095_o = n2094_o;
      4'b0010: n2095_o = n2094_o;
      4'b0001: n2095_o = n2008_o;
      default: n2095_o = n2094_o;
    endcase
  assign n2096_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2097_o = n2096_o;
      4'b0100: n2097_o = n2096_o;
      4'b0010: n2097_o = n2096_o;
      4'b0001: n2097_o = n2019_o;
      default: n2097_o = n2096_o;
    endcase
  assign n2098_o = n1870_o[50];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2099_o = n2098_o;
      4'b0100: n2099_o = n2098_o;
      4'b0010: n2099_o = n2098_o;
      4'b0001: n2099_o = n2017_o;
      default: n2099_o = n2098_o;
    endcase
  assign n2100_o = n1870_o[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2101_o = n2100_o;
      4'b0100: n2101_o = n2100_o;
      4'b0010: n2101_o = n2100_o;
      4'b0001: n2101_o = 1'b1;
      default: n2101_o = n2100_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2102_o = n2071_o;
      4'b0100: n2102_o = n1991_o;
      4'b0010: n2102_o = n1991_o;
      4'b0001: n2102_o = n1991_o;
      default: n2102_o = n1991_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1587:25  */
  always @*
    case (n2079_o)
      4'b1000: n2105_o = n2076_o;
      4'b0100: n2105_o = 7'b0000101;
      4'b0010: n2105_o = 7'b0000100;
      4'b0001: n2105_o = n1968_o;
      default: n2105_o = n1968_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2107_o = n1996_o ? n2082_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2110_o = n1996_o ? n2085_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2113_o = n1996_o ? n2087_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2116_o = n1996_o ? n2089_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2119_o = n1996_o ? n2091_o : 1'b0;
  assign n2121_o = {n2097_o, n2095_o};
  assign n2122_o = n1870_o[22];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2123_o = n1996_o ? n2093_o : n2122_o;
  assign n2124_o = n1870_o[47:46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2125_o = n1996_o ? n2121_o : n2124_o;
  assign n2126_o = n1870_o[50];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2127_o = n1996_o ? n2099_o : n2126_o;
  assign n2128_o = n1870_o[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2129_o = n1996_o ? n2101_o : n2128_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2130_o = n1996_o ? n2102_o : n1991_o;
  assign n2136_o = n1870_o[49:48];
  assign n2137_o = n1870_o[64:63];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n2139_o = n1996_o ? n2105_o : n1968_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:28  */
  assign n2140_o = opcode[15:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:34  */
  assign n2141_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:52  */
  assign n2142_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:64  */
  assign n2144_o = n2142_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:42  */
  assign n2145_o = n2141_o & n2144_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1647:42  */
  assign n2148_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1647:45  */
  assign n2149_o = ~n2148_o;
  assign n2153_o = n1870_o[37];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1647:33  */
  assign n2154_o = n2149_o ? 1'b1 : n2153_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1647:33  */
  assign n2156_o = n2149_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1647:33  */
  assign n2158_o = n2149_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1653:50  */
  assign n2159_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1652:33  */
  assign n2161_o = n2167_o ? 1'b1 : n2154_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1656:50  */
  assign n2162_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1656:53  */
  assign n2163_o = ~n2162_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1652:33  */
  assign n2165_o = n2166_o ? 1'b1 : n2113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1652:33  */
  assign n2166_o = decodeopc & n2163_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1652:33  */
  assign n2167_o = decodeopc & n2159_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1652:33  */
  assign n2169_o = decodeopc ? 7'b1001010 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1661:33  */
  assign n2172_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:42  */
  assign n2173_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:59  */
  assign n2174_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:72  */
  assign n2176_o = n2174_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:50  */
  assign n2177_o = n2173_o | n2176_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:50  */
  assign n2178_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:62  */
  assign n2180_o = n2178_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1667:51  */
  assign n2181_o = opcode[8:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1667:63  */
  assign n2183_o = n2181_o != 6'b000111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1667:83  */
  assign n2184_o = opcode[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1667:86  */
  assign n2185_o = ~n2184_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1667:74  */
  assign n2186_o = n2183_o | n2185_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:70  */
  assign n2187_o = n2180_o & n2186_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1668:51  */
  assign n2188_o = opcode[8:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1668:63  */
  assign n2190_o = n2188_o != 7'b1001111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1668:84  */
  assign n2191_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1668:96  */
  assign n2193_o = n2191_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1668:75  */
  assign n2194_o = n2190_o | n2193_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1667:92  */
  assign n2195_o = n2187_o & n2194_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:51  */
  assign n2196_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:63  */
  assign n2198_o = n2196_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:78  */
  assign n2199_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:90  */
  assign n2201_o = n2199_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:69  */
  assign n2202_o = n2198_o | n2201_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:107  */
  assign n2203_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:119  */
  assign n2205_o = n2203_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1669:98  */
  assign n2206_o = n2202_o | n2205_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1668:103  */
  assign n2207_o = n2195_o & n2206_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1672:58  */
  assign n2210_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1672:70  */
  assign n2212_o = n2210_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1673:66  */
  assign n2213_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1673:78  */
  assign n2215_o = n2213_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1673:57  */
  assign n2218_o = n2215_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1672:49  */
  assign n2221_o = n2212_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1672:49  */
  assign n2223_o = n2212_o ? n2218_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1678:58  */
  assign n2224_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1678:70  */
  assign n2226_o = n2224_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1678:49  */
  assign n2229_o = n2226_o ? 2'b10 : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1683:58  */
  assign n2230_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1683:61  */
  assign n2231_o = ~n2230_o;
  assign n2234_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2235_o = n2260_o ? 1'b1 : n2234_o;
  assign n2236_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2237_o = n2262_o ? 1'b1 : n2236_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2239_o = n2269_o ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1683:49  */
  assign n2242_o = n2231_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1683:49  */
  assign n2244_o = n2231_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1683:49  */
  assign n2246_o = n2231_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1683:49  */
  assign n2247_o = n2231_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2248_o = n2207_o ? n2229_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2250_o = n2207_o ? n2221_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2253_o = n2207_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2256_o = n2207_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2258_o = n2207_o ? n2242_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2260_o = n2207_o & n2244_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2262_o = n2207_o & n2246_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2264_o = n2207_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2266_o = n2207_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2268_o = n2207_o ? n2223_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1666:41  */
  assign n2269_o = n2207_o & n2247_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:45  */
  assign n2270_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:57  */
  assign n2272_o = n2270_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:47  */
  assign n2273_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:58  */
  assign n2274_o = opcode[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:67  */
  assign n2275_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:80  */
  assign n2277_o = n2275_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:66  */
  assign n2278_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:78  */
  assign n2280_o = n2278_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:87  */
  assign n2281_o = n2277_o & n2280_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:96  */
  assign n2282_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:108  */
  assign n2284_o = n2282_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:125  */
  assign n2285_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:137  */
  assign n2287_o = n2285_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:116  */
  assign n2288_o = n2284_o | n2287_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:85  */
  assign n2289_o = n2281_o & n2288_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1701:67  */
  assign n2290_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1701:86  */
  assign n2291_o = opcode[5:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1701:98  */
  assign n2293_o = n2291_o == 6'b111100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1701:76  */
  assign n2294_o = n2290_o & n2293_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1700:145  */
  assign n2295_o = n2289_o | n2294_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1702:76  */
  assign n2296_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1703:73  */
  assign n2298_o = n2296_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1704:73  */
  assign n2300_o = n2296_o == 2'b10;
  assign n2301_o = {n2300_o, n2298_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1702:65  */
  always @*
    case (n2301_o)
      2'b10: n2305_o = 2'b01;
      2'b01: n2305_o = 2'b00;
      default: n2305_o = 2'b10;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:74  */
  assign n2306_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:93  */
  assign n2307_o = opcode[5:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:105  */
  assign n2309_o = n2307_o == 6'b111100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:83  */
  assign n2310_o = n2306_o & n2309_o;
  assign n2312_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1708:73  */
  assign n2313_o = decodeopc ? 1'b1 : n2312_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1708:73  */
  assign n2315_o = decodeopc ? 7'b0111001 : n2139_o;
  assign n2318_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1713:73  */
  assign n2319_o = decodeopc ? 1'b1 : n2318_o;
  assign n2320_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1713:73  */
  assign n2321_o = decodeopc ? 1'b1 : n2320_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1713:73  */
  assign n2323_o = decodeopc ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:87  */
  assign n2325_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:93  */
  assign n2326_o = n2325_o & nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:73  */
  assign n2332_o = n2326_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:73  */
  assign n2335_o = n2326_o ? 1'b1 : 1'b0;
  assign n2336_o = n1870_o[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:73  */
  assign n2337_o = n2326_o ? 1'b1 : n2336_o;
  assign n2338_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:73  */
  assign n2339_o = n2326_o ? 1'b1 : n2338_o;
  assign n2340_o = n1870_o[84];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:73  */
  assign n2341_o = n2326_o ? 1'b1 : n2340_o;
  assign n2342_o = n1870_o[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:73  */
  assign n2343_o = n2326_o ? 1'b1 : n2342_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1718:73  */
  assign n2345_o = n2326_o ? 7'b0110111 : n2323_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2346_o = n2310_o ? n1985_o : n2332_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2348_o = n2310_o ? 1'b0 : n2335_o;
  assign n2349_o = n1870_o[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2350_o = n2310_o ? n2349_o : n2337_o;
  assign n2351_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2352_o = n2310_o ? n2351_o : n2319_o;
  assign n2353_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2354_o = n2310_o ? n2353_o : n2339_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2355_o = n2310_o ? n2313_o : n2321_o;
  assign n2356_o = n1870_o[84];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2357_o = n2310_o ? n2356_o : n2341_o;
  assign n2358_o = n1870_o[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2359_o = n2310_o ? n2358_o : n2343_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1707:65  */
  assign n2360_o = n2310_o ? n2315_o : n2345_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2361_o = n2295_o ? n2305_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2362_o = n2295_o ? n2346_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2364_o = n2295_o ? n2348_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2367_o = n2295_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2370_o = n2295_o ? 1'b0 : 1'b1;
  assign n2371_o = n1870_o[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2372_o = n2950_o ? n2350_o : n2371_o;
  assign n2373_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2374_o = n2295_o ? n2352_o : n2373_o;
  assign n2375_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2376_o = n2479_o ? n2354_o : n2375_o;
  assign n2377_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2378_o = n2295_o ? n2355_o : n2377_o;
  assign n2379_o = n1870_o[84];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2380_o = n2972_o ? n2357_o : n2379_o;
  assign n2381_o = n1870_o[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2382_o = n2974_o ? n2359_o : n2381_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1699:57  */
  assign n2383_o = n2295_o ? n2360_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:66  */
  assign n2384_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:79  */
  assign n2386_o = n2384_o != 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:66  */
  assign n2387_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:78  */
  assign n2389_o = n2387_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:86  */
  assign n2390_o = n2386_o & n2389_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:95  */
  assign n2391_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:107  */
  assign n2393_o = n2391_o != 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:85  */
  assign n2394_o = n2390_o & n2393_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:125  */
  assign n2395_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:137  */
  assign n2397_o = n2395_o != 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:115  */
  assign n2398_o = n2394_o & n2397_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:155  */
  assign n2399_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:167  */
  assign n2401_o = n2399_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1734:145  */
  assign n2402_o = n2398_o & n2401_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1736:83  */
  assign n2404_o = opcode[10:9];
  assign n2407_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1737:65  */
  assign n2408_o = decodeopc ? 1'b1 : n2407_o;
  assign n2409_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2410_o = n2455_o ? 1'b1 : n2409_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1737:65  */
  assign n2412_o = decodeopc ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1742:71  */
  assign n2413_o = set[62];
  assign n2416_o = n1870_o[39];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2417_o = n2449_o ? 1'b1 : n2416_o;
  assign n2418_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2419_o = n2453_o ? 1'b1 : n2418_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1746:79  */
  assign n2421_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1746:85  */
  assign n2422_o = n2421_o & nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1749:88  */
  assign n2425_o = exe_datatype != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1749:73  */
  assign n2428_o = n2425_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2430_o = n2438_o ? 2'b10 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1746:65  */
  assign n2432_o = n2422_o ? n2428_o : 1'b0;
  assign n2433_o = n1870_o[82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2434_o = n2457_o ? 1'b1 : n2433_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1746:65  */
  assign n2436_o = n2422_o ? 7'b1000001 : n2412_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2437_o = n2402_o ? n2404_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2438_o = n2402_o & n2422_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2441_o = n2402_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2444_o = n2402_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2446_o = n2402_o ? n2432_o : 1'b0;
  assign n2447_o = {1'b1, n2408_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2449_o = n2402_o & n2413_o;
  assign n2450_o = n1870_o[43:42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2451_o = n2402_o ? n2447_o : n2450_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2453_o = n2402_o & n2413_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2455_o = n2402_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2457_o = n2402_o & n2422_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1733:57  */
  assign n2458_o = n2402_o ? n2436_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2459_o = n2274_o ? n2361_o : n2437_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2460_o = n2274_o ? n2362_o : n2430_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2462_o = n2274_o ? n2364_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2463_o = n2274_o ? n2367_o : n2441_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2464_o = n2274_o ? n2370_o : n2444_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2466_o = n2274_o ? 1'b0 : n2446_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2468_o = n2274_o & n2295_o;
  assign n2469_o = n1870_o[39];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2470_o = n2274_o ? n2469_o : n2417_o;
  assign n2471_o = n2451_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2472_o = n2274_o ? n2374_o : n2471_o;
  assign n2473_o = n2451_o[1];
  assign n2474_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2475_o = n2274_o ? n2474_o : n2473_o;
  assign n2476_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2477_o = n2274_o ? n2476_o : n2419_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2479_o = n2274_o & n2295_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2480_o = n2274_o ? n2378_o : n2410_o;
  assign n2481_o = n1870_o[82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2482_o = n2274_o ? n2481_o : n2434_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2484_o = n2274_o & n2295_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2486_o = n2274_o & n2295_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1698:49  */
  assign n2487_o = n2274_o ? n2383_o : n2458_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2488_o = n2934_o ? n2459_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2489_o = n2273_o ? n2460_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2491_o = n2273_o ? n2462_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2493_o = n2273_o ? n2463_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2495_o = n2273_o ? n2464_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2497_o = n2273_o ? n2466_o : 1'b0;
  assign n2498_o = {n2475_o, n2472_o};
  assign n2499_o = {n2376_o, n2477_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2501_o = n2273_o & n2468_o;
  assign n2502_o = n1870_o[39];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2503_o = n2952_o ? n2470_o : n2502_o;
  assign n2504_o = n1870_o[43:42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2505_o = n2273_o ? n2498_o : n2504_o;
  assign n2506_o = n1870_o[56:55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2507_o = n2273_o ? n2499_o : n2506_o;
  assign n2508_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2509_o = n2273_o ? n2480_o : n2508_o;
  assign n2510_o = n1870_o[82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2511_o = n2970_o ? n2482_o : n2510_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2513_o = n2273_o & n2484_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2515_o = n2273_o & n2486_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1697:41  */
  assign n2516_o = n2273_o ? n2487_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:45  */
  assign n2517_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:58  */
  assign n2519_o = n2517_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:47  */
  assign n2520_o = cpu[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:65  */
  assign n2521_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:77  */
  assign n2523_o = n2521_o != 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:55  */
  assign n2524_o = n2520_o & n2523_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:94  */
  assign n2525_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:106  */
  assign n2527_o = n2525_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:84  */
  assign n2528_o = n2524_o & n2527_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:124  */
  assign n2529_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:136  */
  assign n2531_o = n2529_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:153  */
  assign n2532_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:165  */
  assign n2534_o = n2532_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:144  */
  assign n2535_o = n2531_o | n2534_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:113  */
  assign n2536_o = n2528_o & n2535_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1765:49  */
  assign n2539_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1765:49  */
  assign n2542_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:41  */
  assign n2544_o = n2536_o ? n2539_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1764:41  */
  assign n2546_o = n2536_o ? n2542_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:50  */
  assign n2547_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:62  */
  assign n2549_o = n2547_o != 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:79  */
  assign n2550_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:91  */
  assign n2552_o = n2550_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:69  */
  assign n2553_o = n2549_o & n2552_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1779:58  */
  assign n2554_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1779:71  */
  assign n2556_o = n2554_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:66  */
  assign n2557_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:78  */
  assign n2559_o = n2557_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:95  */
  assign n2560_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:107  */
  assign n2562_o = n2560_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:86  */
  assign n2563_o = n2559_o | n2562_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:123  */
  assign n2564_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:135  */
  assign n2566_o = n2564_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:152  */
  assign n2567_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:155  */
  assign n2568_o = ~n2567_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:142  */
  assign n2569_o = n2566_o & n2568_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:113  */
  assign n2570_o = n2563_o | n2569_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:57  */
  assign n2574_o = n2570_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:57  */
  assign n2577_o = n2570_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1780:57  */
  assign n2579_o = n2570_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1779:49  */
  assign n2581_o = n2556_o ? n2574_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1779:49  */
  assign n2583_o = n2556_o ? n2577_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1779:49  */
  assign n2585_o = n2556_o ? n2579_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1787:58  */
  assign n2586_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1787:71  */
  assign n2588_o = n2586_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:66  */
  assign n2589_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:78  */
  assign n2591_o = n2589_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:95  */
  assign n2592_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:107  */
  assign n2594_o = n2592_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:86  */
  assign n2595_o = n2591_o | n2594_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:123  */
  assign n2596_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:135  */
  assign n2598_o = n2596_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:152  */
  assign n2599_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:155  */
  assign n2600_o = ~n2599_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:142  */
  assign n2601_o = n2598_o & n2600_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:113  */
  assign n2602_o = n2595_o | n2601_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:57  */
  assign n2605_o = n2602_o ? n2581_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:57  */
  assign n2607_o = n2602_o ? n2583_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1788:57  */
  assign n2609_o = n2602_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1787:49  */
  assign n2610_o = n2588_o ? n2605_o : n2581_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1787:49  */
  assign n2611_o = n2588_o ? n2607_o : n2583_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1787:49  */
  assign n2613_o = n2588_o ? n2609_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:58  */
  assign n2614_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:71  */
  assign n2616_o = n2614_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:87  */
  assign n2617_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:100  */
  assign n2619_o = n2617_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:78  */
  assign n2620_o = n2616_o | n2619_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:66  */
  assign n2621_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:78  */
  assign n2623_o = n2621_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:95  */
  assign n2624_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:107  */
  assign n2626_o = n2624_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:86  */
  assign n2627_o = n2623_o | n2626_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:57  */
  assign n2630_o = n2627_o ? n2610_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:57  */
  assign n2632_o = n2627_o ? n2611_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1796:57  */
  assign n2634_o = n2627_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:49  */
  assign n2635_o = n2620_o ? n2630_o : n2610_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:49  */
  assign n2636_o = n2620_o ? n2632_o : n2611_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1795:49  */
  assign n2638_o = n2620_o ? n2634_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1803:58  */
  assign n2639_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1803:71  */
  assign n2641_o = n2639_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:66  */
  assign n2642_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:78  */
  assign n2644_o = n2642_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:95  */
  assign n2645_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:107  */
  assign n2647_o = n2645_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:86  */
  assign n2648_o = n2644_o | n2647_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:123  */
  assign n2649_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:135  */
  assign n2651_o = n2649_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:152  */
  assign n2652_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:155  */
  assign n2653_o = ~n2652_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:142  */
  assign n2654_o = n2651_o & n2653_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:113  */
  assign n2655_o = n2648_o | n2654_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:57  */
  assign n2658_o = n2655_o ? n2635_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:57  */
  assign n2660_o = n2655_o ? n2636_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1804:57  */
  assign n2662_o = n2655_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1803:49  */
  assign n2663_o = n2641_o ? n2658_o : n2635_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1803:49  */
  assign n2664_o = n2641_o ? n2660_o : n2636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1803:49  */
  assign n2666_o = n2641_o ? n2662_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1811:58  */
  assign n2667_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1811:71  */
  assign n2669_o = n2667_o == 3'b110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:66  */
  assign n2670_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:78  */
  assign n2672_o = n2670_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:95  */
  assign n2673_o = opcode[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:98  */
  assign n2674_o = ~n2673_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:86  */
  assign n2675_o = n2672_o | n2674_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:57  */
  assign n2678_o = n2675_o ? n2663_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:57  */
  assign n2680_o = n2675_o ? n2664_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1812:57  */
  assign n2682_o = n2675_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1811:49  */
  assign n2683_o = n2669_o ? n2678_o : n2663_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1811:49  */
  assign n2684_o = n2669_o ? n2680_o : n2664_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1811:49  */
  assign n2686_o = n2669_o ? n2682_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:61  */
  assign n2687_o = set_exec[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:80  */
  assign n2688_o = set_exec[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:69  */
  assign n2689_o = n2687_o | n2688_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:100  */
  assign n2690_o = set_exec[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:89  */
  assign n2691_o = n2689_o | n2690_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:120  */
  assign n2692_o = set_exec[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:109  */
  assign n2693_o = n2691_o | n2692_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:140  */
  assign n2694_o = set_exec[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:129  */
  assign n2695_o = n2693_o | n2694_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:66  */
  assign n2696_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:69  */
  assign n2697_o = ~n2696_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:84  */
  assign n2698_o = opcode[5:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:96  */
  assign n2700_o = n2698_o == 6'b111100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:74  */
  assign n2701_o = n2697_o & n2700_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:119  */
  assign n2702_o = set_exec[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:139  */
  assign n2703_o = set_exec[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:128  */
  assign n2704_o = n2702_o | n2703_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:158  */
  assign n2705_o = set_exec[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:147  */
  assign n2706_o = n2704_o | n2705_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:106  */
  assign n2707_o = n2701_o & n2706_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:92  */
  assign n2708_o = ~svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:82  */
  assign n2709_o = decodeopc & n2708_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:107  */
  assign n2710_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:97  */
  assign n2711_o = n2709_o & n2710_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1827:90  */
  assign n2713_o = opcode[6];
  assign n2715_o = n1870_o[52];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1827:81  */
  assign n2716_o = n2713_o ? 1'b1 : n2715_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1831:104  */
  assign n2718_o = set_exec[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1832:104  */
  assign n2719_o = set_exec[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1833:103  */
  assign n2720_o = set_exec[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1826:73  */
  assign n2722_o = decodeopc ? 2'b01 : n1985_o;
  assign n2723_o = {n2720_o, n2719_o, n2718_o};
  assign n2724_o = {n2716_o, 1'b1};
  assign n2725_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1826:73  */
  assign n2726_o = decodeopc ? n2723_o : n2725_o;
  assign n2727_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1826:73  */
  assign n2728_o = decodeopc ? n2724_o : n2727_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1826:73  */
  assign n2730_o = decodeopc ? 7'b0011000 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:65  */
  assign n2731_o = n2711_o ? n1985_o : n2722_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:65  */
  assign n2734_o = n2711_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:65  */
  assign n2736_o = n2711_o ? 1'b1 : n2684_o;
  assign n2737_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:65  */
  assign n2738_o = n2711_o ? n2737_o : n2726_o;
  assign n2739_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:65  */
  assign n2740_o = n2711_o ? n2739_o : 1'b1;
  assign n2741_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:65  */
  assign n2742_o = n2711_o ? n2741_o : n2728_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1821:65  */
  assign n2743_o = n2711_o ? n2139_o : n2730_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:69  */
  assign n2744_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:72  */
  assign n2745_o = ~n2744_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:86  */
  assign n2746_o = opcode[5:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:98  */
  assign n2748_o = n2746_o != 6'b111100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:77  */
  assign n2749_o = n2745_o | n2748_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:121  */
  assign n2750_o = set_exec[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:141  */
  assign n2751_o = set_exec[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:130  */
  assign n2752_o = n2750_o | n2751_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:160  */
  assign n2753_o = set_exec[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:149  */
  assign n2754_o = n2752_o | n2753_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:169  */
  assign n2755_o = ~n2754_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:109  */
  assign n2756_o = n2749_o | n2755_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1844:84  */
  assign n2760_o = datatype == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2762_o = n2811_o ? 1'b1 : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2764_o = n2800_o ? 1'b1 : n2113_o;
  assign n2765_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2766_o = n2806_o ? 1'b1 : n2765_o;
  assign n2767_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2768_o = n2810_o ? 1'b1 : n2767_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1839:65  */
  assign n2769_o = decodeopc & n2760_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2771_o = n2816_o ? 7'b0011101 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1848:74  */
  assign n2772_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1848:86  */
  assign n2774_o = n2772_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1848:65  */
  assign n2777_o = n2774_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1851:74  */
  assign n2778_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1851:87  */
  assign n2780_o = n2778_o != 3'b110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1852:82  */
  assign n2781_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1852:94  */
  assign n2783_o = n2781_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1852:73  */
  assign n2786_o = n2783_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1851:65  */
  assign n2789_o = n2780_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1851:65  */
  assign n2791_o = n2780_o ? n2786_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1857:74  */
  assign n2792_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1857:87  */
  assign n2794_o = n2792_o == 2'b10;
  assign n2796_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2797_o = n2808_o ? 1'b1 : n2796_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2799_o = n2756_o ? n2789_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2800_o = n2756_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2802_o = n2756_o ? n2683_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2804_o = n2756_o ? n2684_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2806_o = n2756_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2808_o = n2756_o & n2794_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2810_o = n2756_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2811_o = n2756_o & n2769_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2813_o = n2756_o ? n2777_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2815_o = n2756_o ? n2791_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1838:57  */
  assign n2816_o = n2756_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2817_o = n2871_o ? n2731_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2819_o = n2707_o ? 1'b0 : n2799_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2820_o = n2707_o ? n2113_o : n2764_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2821_o = n2707_o ? n2683_o : n2802_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2823_o = n2707_o ? n2734_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2824_o = n2707_o ? n2736_o : n2804_o;
  assign n2825_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2826_o = n2882_o ? n2738_o : n2825_o;
  assign n2827_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2828_o = n2707_o ? n2827_o : n2766_o;
  assign n2829_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2830_o = n2886_o ? n2740_o : n2829_o;
  assign n2831_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2832_o = n2888_o ? n2742_o : n2831_o;
  assign n2833_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2834_o = n2707_o ? n2833_o : n2797_o;
  assign n2835_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2836_o = n2707_o ? n2835_o : n2768_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2837_o = n2707_o ? n2130_o : n2762_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2839_o = n2707_o ? 1'b0 : n2813_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2841_o = n2707_o ? 1'b0 : n2815_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1820:57  */
  assign n2842_o = n2707_o ? n2743_o : n2771_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2843_o = n2695_o & n2707_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2845_o = n2695_o ? n2819_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2846_o = n2874_o ? n2820_o : n2113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2848_o = n2695_o ? n2821_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2850_o = n2695_o ? n2823_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2852_o = n2695_o ? n2824_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2854_o = n2695_o & n2707_o;
  assign n2855_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2856_o = n2884_o ? n2828_o : n2855_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2858_o = n2695_o & n2707_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2860_o = n2695_o & n2707_o;
  assign n2861_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2862_o = n2890_o ? n2834_o : n2861_o;
  assign n2863_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2864_o = n2892_o ? n2836_o : n2863_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2865_o = n2893_o ? n2837_o : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2867_o = n2695_o ? n2839_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1819:49  */
  assign n2869_o = n2695_o ? n2841_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2870_o = n2903_o ? n2842_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2871_o = n2553_o & n2843_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2873_o = n2553_o ? n2845_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2874_o = n2553_o & n2695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2876_o = n2553_o ? n2848_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2878_o = n2553_o ? n2850_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2880_o = n2553_o ? n2852_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2882_o = n2553_o & n2854_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2884_o = n2553_o & n2695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2886_o = n2553_o & n2858_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2888_o = n2553_o & n2860_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2890_o = n2553_o & n2695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2892_o = n2553_o & n2695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2893_o = n2553_o & n2695_o;
  assign n2894_o = {n2686_o, n2666_o, n2613_o, n2585_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2896_o = n2553_o ? n2638_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2898_o = n2553_o ? n2894_o : 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2900_o = n2553_o ? n2867_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2902_o = n2553_o ? n2869_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1778:41  */
  assign n2903_o = n2553_o & n2695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2904_o = n2519_o ? n1985_o : n2817_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2906_o = n2519_o ? 1'b0 : n2873_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2907_o = n2519_o ? n2113_o : n2846_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2908_o = n2519_o ? n2544_o : n2876_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2909_o = n2519_o ? n2546_o : n2878_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2911_o = n2519_o ? 1'b1 : n2880_o;
  assign n2912_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2913_o = n2519_o ? n2912_o : n2826_o;
  assign n2914_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2915_o = n2519_o ? n2914_o : n2856_o;
  assign n2916_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2917_o = n2519_o ? n2916_o : n2830_o;
  assign n2918_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2919_o = n2519_o ? n2918_o : n2832_o;
  assign n2920_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2921_o = n2519_o ? n2920_o : n2862_o;
  assign n2922_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2923_o = n2519_o ? n2922_o : n2864_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2924_o = n2519_o ? n2130_o : n2865_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2926_o = n2519_o ? 1'b0 : n2896_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2928_o = n2519_o ? 4'b0000 : n2898_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2930_o = n2519_o ? 1'b0 : n2900_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2932_o = n2519_o ? 1'b0 : n2902_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1763:33  */
  assign n2933_o = n2519_o ? n2139_o : n2870_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2934_o = n2272_o & n2273_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2935_o = n2272_o ? n2489_o : n2904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2937_o = n2272_o ? 1'b0 : n2906_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2939_o = n2272_o ? n2491_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2940_o = n2272_o ? n2113_o : n2907_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2941_o = n2272_o ? n2493_o : n2908_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2943_o = n2272_o ? 1'b0 : n2909_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2944_o = n2272_o ? n2495_o : n2911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2946_o = n2272_o ? n2497_o : 1'b0;
  assign n2947_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2948_o = n2272_o ? n2947_o : n2913_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2950_o = n2272_o & n2501_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2952_o = n2272_o & n2273_o;
  assign n2953_o = n2505_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2954_o = n2272_o ? n2953_o : n2915_o;
  assign n2955_o = n2505_o[1];
  assign n2956_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2957_o = n2272_o ? n2955_o : n2956_o;
  assign n2958_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2959_o = n2272_o ? n2958_o : n2917_o;
  assign n2960_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2961_o = n2272_o ? n2960_o : n2919_o;
  assign n2962_o = n2507_o[0];
  assign n2963_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2964_o = n2272_o ? n2962_o : n2963_o;
  assign n2965_o = n2507_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2966_o = n2272_o ? n2965_o : n2921_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2967_o = n2272_o ? n2509_o : n2923_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2968_o = n2272_o ? n2130_o : n2924_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2970_o = n2272_o & n2273_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2972_o = n2272_o & n2513_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2974_o = n2272_o & n2515_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2976_o = n2272_o ? 1'b0 : n2926_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2978_o = n2272_o ? 4'b0000 : n2928_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2980_o = n2272_o ? 1'b0 : n2930_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2982_o = n2272_o ? 1'b0 : n2932_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1696:33  */
  assign n2983_o = n2272_o ? n2516_o : n2933_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2984_o = n2177_o ? n2248_o : n2488_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2985_o = n2177_o ? n1985_o : n2935_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2986_o = n2177_o ? n2250_o : n2937_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2988_o = n2177_o ? 1'b0 : n2939_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2989_o = n2177_o ? n2113_o : n2940_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2990_o = n2177_o ? n2253_o : n2941_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2992_o = n2177_o ? 1'b0 : n2943_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2993_o = n2177_o ? n2256_o : n2944_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2995_o = n2177_o ? n2258_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n2997_o = n2177_o ? 1'b0 : n2946_o;
  assign n2998_o = {n2957_o, n2954_o};
  assign n2999_o = {n2966_o, n2964_o};
  assign n3000_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3001_o = n2177_o ? n3000_o : n2948_o;
  assign n3002_o = n1870_o[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3003_o = n2177_o ? n3002_o : n2372_o;
  assign n3004_o = n1870_o[39];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3005_o = n2177_o ? n3004_o : n2503_o;
  assign n3006_o = n2998_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3007_o = n2177_o ? n2235_o : n3006_o;
  assign n3008_o = n2998_o[1];
  assign n3009_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3010_o = n2177_o ? n3009_o : n3008_o;
  assign n3011_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3012_o = n2177_o ? n3011_o : n2959_o;
  assign n3013_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3014_o = n2177_o ? n3013_o : n2961_o;
  assign n3015_o = n1870_o[56:55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3016_o = n2177_o ? n3015_o : n2999_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3017_o = n2177_o ? n2237_o : n2967_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3018_o = n2177_o ? n2130_o : n2968_o;
  assign n3019_o = n1870_o[82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3020_o = n2177_o ? n3019_o : n2511_o;
  assign n3021_o = n1870_o[84];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3022_o = n2177_o ? n3021_o : n2380_o;
  assign n3023_o = n1870_o[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3024_o = n2177_o ? n3023_o : n2382_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3026_o = n2177_o ? 1'b0 : n2976_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3028_o = n2177_o ? 4'b0000 : n2978_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3030_o = n2177_o ? n2264_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3031_o = n2177_o ? n2266_o : n2980_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3032_o = n2177_o ? n2268_o : n2982_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1665:33  */
  assign n3033_o = n2177_o ? n2239_o : n2983_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3035_o = n2145_o ? 2'b00 : n2984_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3036_o = n2145_o ? n1985_o : n2985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3038_o = n2145_o ? 1'b0 : n2986_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3040_o = n2145_o ? 1'b0 : n2988_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3042_o = n2145_o ? n2172_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3043_o = n2145_o ? n2165_o : n2989_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3045_o = n2145_o ? 1'b0 : n2990_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3047_o = n2145_o ? 1'b0 : n2992_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3049_o = n2145_o ? 1'b0 : n2993_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3051_o = n2145_o ? 1'b0 : n2995_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3053_o = n2145_o ? 1'b0 : n2997_o;
  assign n3054_o = {n3010_o, n3007_o};
  assign n3055_o = {1'b1, 1'b1};
  assign n3056_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3057_o = n2145_o ? n3056_o : n3001_o;
  assign n3058_o = n1870_o[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3059_o = n2145_o ? n3058_o : n3003_o;
  assign n3060_o = n1870_o[37];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3061_o = n2145_o ? n2161_o : n3060_o;
  assign n3062_o = n1870_o[39];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3063_o = n2145_o ? n3062_o : n3005_o;
  assign n3064_o = n1870_o[43:42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3065_o = n2145_o ? n3064_o : n3054_o;
  assign n3066_o = n3055_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3067_o = n2145_o ? n3066_o : n3012_o;
  assign n3068_o = n3055_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3069_o = n2145_o ? n3068_o : n2127_o;
  assign n3070_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3071_o = n2145_o ? n3070_o : n3014_o;
  assign n3072_o = n1870_o[56:55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3073_o = n2145_o ? n3072_o : n3016_o;
  assign n3074_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3075_o = n2145_o ? n3074_o : n3017_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3076_o = n2145_o ? n2130_o : n3018_o;
  assign n3077_o = n1870_o[82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3078_o = n2145_o ? n3077_o : n3020_o;
  assign n3079_o = n1870_o[84];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3080_o = n2145_o ? n3079_o : n3022_o;
  assign n3081_o = n1870_o[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3082_o = n2145_o ? n3081_o : n3024_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3084_o = n2145_o ? n2156_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3086_o = n2145_o ? 1'b0 : n3026_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3088_o = n2145_o ? 4'b0000 : n3028_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3090_o = n2145_o ? 1'b0 : n3030_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3092_o = n2145_o ? 1'b0 : n3031_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3093_o = n2145_o ? n2158_o : n3032_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1643:25  */
  assign n3094_o = n2145_o ? n2169_o : n3033_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1642:25  */
  assign n3096_o = n2140_o == 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:44  */
  assign n3097_o = opcode[11:10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:58  */
  assign n3099_o = n3097_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:73  */
  assign n3100_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:85  */
  assign n3102_o = n3100_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:64  */
  assign n3103_o = n3099_o | n3102_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1878:43  */
  assign n3104_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1878:55  */
  assign n3106_o = n3104_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1878:73  */
  assign n3107_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1878:85  */
  assign n3109_o = n3107_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1878:64  */
  assign n3110_o = n3106_o | n3109_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:94  */
  assign n3111_o = n3103_o & n3110_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1879:43  */
  assign n3112_o = opcode[13];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1879:62  */
  assign n3113_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1879:74  */
  assign n3115_o = n3113_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1879:92  */
  assign n3116_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1879:104  */
  assign n3118_o = n3116_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1879:82  */
  assign n3119_o = n3115_o & n3118_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1879:52  */
  assign n3120_o = n3112_o | n3119_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1878:92  */
  assign n3121_o = n3111_o & n3120_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1882:50  */
  assign n3123_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1882:62  */
  assign n3125_o = n3123_o == 3'b001;
  assign n3127_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1882:41  */
  assign n3128_o = n3125_o ? 1'b1 : n3127_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1885:50  */
  assign n3129_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1885:62  */
  assign n3131_o = n3129_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1886:58  */
  assign n3132_o = opcode[8:7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1886:70  */
  assign n3134_o = n3132_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1886:49  */
  assign n3137_o = n3134_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1885:41  */
  assign n3139_o = n3131_o ? n3137_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1890:52  */
  assign n3140_o = opcode[13:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1891:49  */
  assign n3142_o = n3140_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1892:49  */
  assign n3144_o = n3140_o == 2'b10;
  assign n3145_o = {n3144_o, n3142_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1890:41  */
  always @*
    case (n3145_o)
      2'b10: n3149_o = 2'b10;
      2'b01: n3149_o = 2'b00;
      default: n3149_o = 2'b01;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1896:50  */
  assign n3150_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1896:41  */
  assign n3153_o = n3150_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1900:66  */
  assign n3154_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1900:78  */
  assign n3156_o = n3154_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1900:57  */
  assign n3157_o = nextpass | n3156_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1902:58  */
  assign n3158_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1902:70  */
  assign n3160_o = n3158_o != 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1902:49  */
  assign n3163_o = n3160_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1900:41  */
  assign n3165_o = n3157_o ? n3163_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1900:41  */
  assign n3168_o = n3157_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:55  */
  assign n3170_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:89  */
  assign n3171_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:101  */
  assign n3173_o = n3171_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:107  */
  assign n3174_o = n3173_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:79  */
  assign n3175_o = nextpass | n3174_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:61  */
  assign n3176_o = n3170_o & n3175_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:60  */
  assign n3177_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1909:57  */
  assign n3180_o = n3177_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1909:67  */
  assign n3182_o = n3177_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1909:67  */
  assign n3183_o = n3180_o | n3182_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1912:74  */
  assign n3184_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1914:82  */
  assign n3186_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1914:95  */
  assign n3188_o = n3186_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1912:65  */
  assign n3190_o = n3195_o ? 1'b1 : n2127_o;
  assign n3191_o = n2121_o[0];
  assign n3192_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n3193_o = n1996_o ? n3191_o : n3192_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1912:65  */
  assign n3194_o = n3184_o ? 1'b1 : n3193_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1912:65  */
  assign n3195_o = n3184_o & n3188_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1918:74  */
  assign n3196_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1920:82  */
  assign n3198_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1920:95  */
  assign n3200_o = n3198_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1918:65  */
  assign n3202_o = n3207_o ? 1'b1 : n3190_o;
  assign n3203_o = n2121_o[1];
  assign n3204_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n3205_o = n1996_o ? n3203_o : n3204_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1918:65  */
  assign n3206_o = n3196_o ? 1'b1 : n3205_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1918:65  */
  assign n3207_o = n3196_o & n3200_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1926:76  */
  assign n3208_o = ~nextpass;
  assign n3210_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1926:65  */
  assign n3211_o = n3208_o ? 1'b1 : n3210_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1911:57  */
  assign n3213_o = n3177_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1911:67  */
  assign n3215_o = n3177_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1911:67  */
  assign n3216_o = n3213_o | n3215_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1911:73  */
  assign n3218_o = n3177_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1911:73  */
  assign n3219_o = n3216_o | n3218_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1929:57  */
  assign n3221_o = n3177_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1932:57  */
  assign n3223_o = n3177_o == 3'b110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1936:76  */
  assign n3224_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1937:73  */
  assign n3226_o = n3224_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1939:73  */
  assign n3229_o = n3224_o == 3'b001;
  assign n3230_o = {n3229_o, n3226_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1936:65  */
  always @*
    case (n3230_o)
      2'b10: n3231_o = 1'b1;
      2'b01: n3231_o = n2130_o;
      default: n3231_o = n2130_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1936:65  */
  always @*
    case (n3230_o)
      2'b10: n3234_o = 7'b0000011;
      2'b01: n3234_o = 7'b0000011;
      default: n3234_o = n2139_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1935:57  */
  assign n3236_o = n3177_o == 3'b111;
  assign n3237_o = {n3236_o, n3223_o, n3221_o, n3219_o, n3183_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3239_o = n1985_o;
      5'b01000: n3239_o = n1985_o;
      5'b00100: n3239_o = n1985_o;
      5'b00010: n3239_o = 2'b11;
      5'b00001: n3239_o = n1985_o;
      default: n3239_o = n1985_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3241_o = n2110_o;
      5'b01000: n3241_o = 1'b1;
      5'b00100: n3241_o = n2110_o;
      5'b00010: n3241_o = n2110_o;
      5'b00001: n3241_o = n2110_o;
      default: n3241_o = n2110_o;
    endcase
  assign n3242_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3243_o = n3242_o;
      5'b01000: n3243_o = n3242_o;
      5'b00100: n3243_o = n3242_o;
      5'b00010: n3243_o = n3211_o;
      5'b00001: n3243_o = n3242_o;
      default: n3243_o = n3242_o;
    endcase
  assign n3244_o = n2121_o[0];
  assign n3245_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n3246_o = n1996_o ? n3244_o : n3245_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3247_o = n3246_o;
      5'b01000: n3247_o = n3246_o;
      5'b00100: n3247_o = n3246_o;
      5'b00010: n3247_o = n3194_o;
      5'b00001: n3247_o = n3246_o;
      default: n3247_o = n3246_o;
    endcase
  assign n3248_o = n2121_o[1];
  assign n3249_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n3250_o = n1996_o ? n3248_o : n3249_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3251_o = n3250_o;
      5'b01000: n3251_o = n3250_o;
      5'b00100: n3251_o = n3250_o;
      5'b00010: n3251_o = n3206_o;
      5'b00001: n3251_o = n3250_o;
      default: n3251_o = n3250_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3252_o = n2127_o;
      5'b01000: n3252_o = n2127_o;
      5'b00100: n3252_o = n2127_o;
      5'b00010: n3252_o = n3202_o;
      5'b00001: n3252_o = n2127_o;
      default: n3252_o = n2127_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3253_o = n3231_o;
      5'b01000: n3253_o = n2130_o;
      5'b00100: n3253_o = n2130_o;
      5'b00010: n3253_o = n2130_o;
      5'b00001: n3253_o = n2130_o;
      default: n3253_o = n2130_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3254_o = n3139_o;
      5'b01000: n3254_o = n3139_o;
      5'b00100: n3254_o = n3139_o;
      5'b00010: n3254_o = n3139_o;
      5'b00001: n3254_o = 1'b1;
      default: n3254_o = n3139_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1908:49  */
  always @*
    case (n3237_o)
      5'b10000: n3258_o = n3234_o;
      5'b01000: n3258_o = 7'b0010011;
      5'b00100: n3258_o = 7'b0000111;
      5'b00010: n3258_o = 7'b0000001;
      5'b00001: n3258_o = n2139_o;
      default: n3258_o = n2139_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3259_o = n3270_o ? n3239_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3260_o = n3271_o ? n3241_o : n2110_o;
  assign n3261_o = {n3251_o, n3247_o};
  assign n3262_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3263_o = n3292_o ? n3243_o : n3262_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3264_o = n3293_o ? n3261_o : n2125_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:41  */
  assign n3265_o = n3176_o ? n3252_o : n2127_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3266_o = n3297_o ? n3253_o : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1907:41  */
  assign n3267_o = n3176_o ? n3254_o : n3139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3268_o = n3302_o ? n3258_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3269_o = n3121_o ? n3149_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3270_o = n3121_o & n3176_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3271_o = n3121_o & n3176_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3273_o = n3121_o ? n3153_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3276_o = n3121_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3278_o = n3121_o ? n3165_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3280_o = n3121_o ? n3168_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3283_o = n3121_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3286_o = n3121_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3289_o = n3121_o ? 1'b1 : 1'b0;
  assign n3290_o = {n3265_o, n3128_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3292_o = n3121_o & n3176_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3293_o = n3121_o & n3176_o;
  assign n3294_o = n1870_o[49];
  assign n3295_o = {n2127_o, n3294_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3296_o = n3121_o ? n3290_o : n3295_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3297_o = n3121_o & n3176_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3299_o = n3121_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3301_o = n3121_o ? n3267_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1877:33  */
  assign n3302_o = n3121_o & n3176_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1876:25  */
  assign n3304_o = n2140_o == 4'b0001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1876:36  */
  assign n3306_o = n2140_o == 4'b0010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1876:36  */
  assign n3307_o = n3304_o | n3306_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1876:43  */
  assign n3309_o = n2140_o == 4'b0011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1876:43  */
  assign n3310_o = n3307_o | n3309_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:42  */
  assign n3311_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:50  */
  assign n3312_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:58  */
  assign n3313_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:71  */
  assign n3315_o = n3313_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:88  */
  assign n3316_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:100  */
  assign n3318_o = n3316_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:78  */
  assign n3319_o = n3315_o & n3318_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:66  */
  assign n3320_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:81  */
  assign n3321_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:74  */
  assign n3322_o = n3320_o & n3321_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:57  */
  assign n3329_o = n3322_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:57  */
  assign n3332_o = n3322_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:57  */
  assign n3335_o = n3322_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:57  */
  assign n3337_o = n3322_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:57  */
  assign n3339_o = n3322_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:57  */
  assign n3341_o = n3322_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1956:57  */
  assign n3343_o = n3322_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:66  */
  assign n3344_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1968:67  */
  assign n3345_o = opcode[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1968:84  */
  assign n3346_o = opcode[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1968:96  */
  assign n3348_o = n3346_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1968:75  */
  assign n3349_o = n3345_o | n3348_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:74  */
  assign n3350_o = n3344_o & n3349_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1969:66  */
  assign n3351_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1969:78  */
  assign n3353_o = n3351_o != 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1968:103  */
  assign n3354_o = n3350_o & n3353_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1969:96  */
  assign n3355_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1969:108  */
  assign n3357_o = n3355_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1969:86  */
  assign n3358_o = n3354_o & n3357_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1976:74  */
  assign n3362_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1976:86  */
  assign n3364_o = n3362_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1976:65  */
  assign n3367_o = n3364_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1976:65  */
  assign n3370_o = n3364_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1976:65  */
  assign n3373_o = n3364_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1982:71  */
  assign n3374_o = set[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3376_o = n3383_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3378_o = n3397_o ? 1'b1 : n2113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1986:65  */
  assign n3380_o = setexecopc ? 1'b1 : n3367_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1986:65  */
  assign n3382_o = setexecopc ? 1'b1 : n3370_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3383_o = n3358_o & n3374_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3386_o = n3358_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3389_o = n3358_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3392_o = n3358_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3394_o = n3358_o ? n3380_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3396_o = n3358_o ? n3382_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3397_o = n3358_o & n3374_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3400_o = n3358_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3403_o = n3358_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3405_o = n3358_o ? n3373_o : 1'b0;
  assign n3406_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3407_o = n3358_o ? 1'b1 : n3406_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3409_o = n3358_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1967:57  */
  assign n3411_o = n3358_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3412_o = n3319_o ? n1985_o : n3376_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3414_o = n3319_o ? 1'b0 : n3386_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3416_o = n3319_o ? 1'b0 : n3389_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3417_o = n3319_o ? n3329_o : n3392_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3419_o = n3319_o ? 1'b0 : n3394_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3421_o = n3319_o ? 1'b0 : n3396_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3422_o = n3319_o ? n2113_o : n3378_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3423_o = n3319_o ? n3332_o : n3400_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3424_o = n3319_o ? n3335_o : n3403_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3426_o = n3319_o ? 1'b0 : n3405_o;
  assign n3427_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3428_o = n3319_o ? n3427_o : n3407_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3429_o = n3319_o ? n3337_o : n3409_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3431_o = n3319_o ? n3339_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3432_o = n3319_o ? n3341_o : n3411_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1955:49  */
  assign n3434_o = n3319_o ? n3343_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:58  */
  assign n3435_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:70  */
  assign n3437_o = n3435_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1997:59  */
  assign n3438_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1997:71  */
  assign n3440_o = n3438_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1997:89  */
  assign n3441_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1997:101  */
  assign n3443_o = n3441_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1997:80  */
  assign n3444_o = n3440_o | n3443_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:78  */
  assign n3445_o = n3437_o & n3444_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1998:66  */
  assign n3446_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:74  */
  assign n3448_o = c_out[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:77  */
  assign n3449_o = ~n3448_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:91  */
  assign n3450_o = op1out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:82  */
  assign n3451_o = n3449_o | n3450_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:109  */
  assign n3452_o = op2out[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:100  */
  assign n3453_o = n3451_o | n3452_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:127  */
  assign n3454_o = exec[31];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:119  */
  assign n3455_o = n3453_o & n3454_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2001:65  */
  assign n3458_o = n3455_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2004:66  */
  assign n3459_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:74  */
  assign n3461_o = c_out[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:77  */
  assign n3462_o = ~n3461_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:91  */
  assign n3463_o = op1out[31];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:82  */
  assign n3464_o = n3462_o | n3463_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:109  */
  assign n3465_o = op2out[31];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:100  */
  assign n3466_o = n3464_o | n3465_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:127  */
  assign n3467_o = exec[31];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:119  */
  assign n3468_o = n3466_o & n3467_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2007:65  */
  assign n3471_o = n3468_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2004:57  */
  assign n3473_o = n3459_o ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2004:57  */
  assign n3476_o = n3459_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2004:57  */
  assign n3478_o = n3459_o ? n3471_o : 1'b1;
  assign n3479_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2004:57  */
  assign n3480_o = n3459_o ? 1'b1 : n3479_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1998:57  */
  assign n3482_o = n3446_o ? 2'b01 : n3473_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1998:57  */
  assign n3484_o = n3446_o ? 1'b0 : n3476_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1998:57  */
  assign n3485_o = n3446_o ? n3458_o : n3478_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1998:57  */
  assign n3486_o = n3446_o ? 1'b1 : n3480_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2014:66  */
  assign n3487_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2014:80  */
  assign n3488_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2014:74  */
  assign n3489_o = n3487_o | n3488_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:91  */
  assign n3490_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:103  */
  assign n3492_o = n3490_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:82  */
  assign n3493_o = nextpass | n3492_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:118  */
  assign n3494_o = exec[31];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:126  */
  assign n3495_o = ~n3494_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:110  */
  assign n3496_o = n3493_o & n3495_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:146  */
  assign n3498_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:131  */
  assign n3499_o = n3496_o & n3498_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2015:65  */
  assign n3502_o = n3499_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2020:65  */
  assign n3506_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2020:65  */
  assign n3509_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2014:57  */
  assign n3511_o = n3489_o ? n3506_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2014:57  */
  assign n3513_o = n3489_o ? n3509_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2014:57  */
  assign n3516_o = n3489_o ? 1'b1 : 1'b0;
  assign n3517_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3518_o = n3535_o ? 1'b1 : n3517_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2014:57  */
  assign n3520_o = n3489_o ? n3502_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3521_o = n3445_o ? n3482_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3523_o = n3445_o ? n3511_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3525_o = n3445_o ? n3513_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3527_o = n3445_o ? n3484_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3529_o = n3445_o ? n3485_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3531_o = n3445_o ? n3516_o : 1'b0;
  assign n3532_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3533_o = n3445_o ? n3486_o : n3532_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3535_o = n3445_o & n3489_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1996:49  */
  assign n3537_o = n3445_o ? n3520_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3538_o = n3312_o ? n1882_o : n3521_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3539_o = n3312_o ? n3412_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3541_o = n3312_o ? n3414_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3543_o = n3312_o ? n3416_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3544_o = n3312_o ? n3417_o : n3523_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3546_o = n3312_o ? n3419_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3547_o = n3312_o ? n3421_o : n3525_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3548_o = n3312_o ? n3422_o : n2113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3549_o = n3312_o ? n3423_o : n3527_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3550_o = n3312_o ? n3424_o : n3529_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3551_o = n3312_o ? n3426_o : n3531_o;
  assign n3552_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3553_o = n3312_o ? n3552_o : n3533_o;
  assign n3554_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3555_o = n3312_o ? n3428_o : n3554_o;
  assign n3556_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3557_o = n3312_o ? n3556_o : n3518_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3559_o = n3312_o ? n3429_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3561_o = n3312_o ? n3431_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3563_o = n3312_o ? 1'b0 : n3537_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3565_o = n3312_o ? n3432_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1954:41  */
  assign n3567_o = n3312_o ? n3434_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:52  */
  assign n3568_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:67  */
  assign n3569_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:79  */
  assign n3571_o = n3569_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2034:67  */
  assign n3572_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2034:79  */
  assign n3574_o = n3572_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2034:96  */
  assign n3575_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2034:108  */
  assign n3577_o = n3575_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2034:87  */
  assign n3578_o = n3574_o | n3577_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:87  */
  assign n3579_o = n3571_o & n3578_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:74  */
  assign n3580_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:86  */
  assign n3582_o = n3580_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:93  */
  assign n3583_o = cpu[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:96  */
  assign n3584_o = ~n3583_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:101  */
  assign n3586_o = n3584_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:86  */
  assign n3588_o = 1'b0 | n3586_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:116  */
  assign n3589_o = n3588_o | svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2041:87  */
  assign n3591_o = cpu[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2041:104  */
  assign n3593_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2041:95  */
  assign n3594_o = n3591_o & n3593_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2041:123  */
  assign n3595_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2041:110  */
  assign n3596_o = n3594_o & n3595_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3598_o = n3660_o ? 1'b1 : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2044:90  */
  assign n3599_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2044:102  */
  assign n3601_o = n3599_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2044:81  */
  assign n3604_o = n3601_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:73  */
  assign n3605_o = n3589_o & n3596_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3607_o = n3661_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:73  */
  assign n3610_o = n3589_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:73  */
  assign n3613_o = n3589_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:73  */
  assign n3616_o = n3589_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:73  */
  assign n3619_o = n3589_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:73  */
  assign n3621_o = n3589_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2036:73  */
  assign n3623_o = n3589_o ? n3604_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2058:82  */
  assign n3627_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2058:94  */
  assign n3629_o = n3627_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2058:73  */
  assign n3632_o = n3629_o ? 1'b1 : 1'b0;
  assign n3634_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2061:73  */
  assign n3635_o = setexecopc ? 1'b1 : n3634_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3636_o = n3582_o & n3605_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3637_o = n3582_o & n3589_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3639_o = n3582_o ? n3610_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3642_o = n3582_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3644_o = n3582_o ? n3613_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3646_o = n3582_o ? n3616_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3648_o = n3582_o ? n3619_o : 1'b1;
  assign n3649_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3650_o = n3582_o ? n3649_o : n3635_o;
  assign n3651_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3652_o = n3582_o ? n3651_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3654_o = n3582_o ? n3621_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3656_o = n3582_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3658_o = n3582_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2035:65  */
  assign n3659_o = n3582_o ? n3623_o : n3632_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3660_o = n3579_o & n3636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3661_o = n3579_o & n3637_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3663_o = n3579_o ? n3639_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3665_o = n3579_o ? n3642_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3668_o = n3579_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3670_o = n3579_o ? n3644_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3672_o = n3579_o ? n3646_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3674_o = n3579_o ? n3648_o : 1'b0;
  assign n3675_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3676_o = n3579_o ? n3650_o : n3675_o;
  assign n3677_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3678_o = n3579_o ? n3652_o : n3677_o;
  assign n3679_o = {n3656_o, n3654_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3681_o = n3579_o ? n3679_o : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3683_o = n3579_o ? n3658_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2033:57  */
  assign n3685_o = n3579_o ? n3659_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2032:49  */
  assign n3687_o = n3568_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:67  */
  assign n3688_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:79  */
  assign n3690_o = n3688_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2071:67  */
  assign n3691_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2071:79  */
  assign n3693_o = n3691_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2071:96  */
  assign n3694_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2071:108  */
  assign n3696_o = n3694_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2071:87  */
  assign n3697_o = n3693_o | n3696_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:87  */
  assign n3698_o = n3690_o & n3697_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:74  */
  assign n3699_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:86  */
  assign n3701_o = n3699_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:93  */
  assign n3702_o = cpu[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:101  */
  assign n3704_o = n3702_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:86  */
  assign n3706_o = 1'b0 | n3704_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2081:90  */
  assign n3708_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2081:102  */
  assign n3710_o = n3708_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2081:81  */
  assign n3713_o = n3710_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3715_o = n3768_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:73  */
  assign n3718_o = n3706_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:73  */
  assign n3721_o = n3706_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:73  */
  assign n3724_o = n3706_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:73  */
  assign n3727_o = n3706_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:73  */
  assign n3729_o = n3706_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2073:73  */
  assign n3731_o = n3706_o ? n3713_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2092:71  */
  assign n3733_o = cpu[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2092:88  */
  assign n3735_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2092:79  */
  assign n3736_o = n3733_o & n3735_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2092:107  */
  assign n3737_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2092:94  */
  assign n3738_o = n3736_o & n3737_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2092:65  */
  assign n3740_o = n3738_o ? 1'b1 : make_berr;
  assign n3742_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2095:73  */
  assign n3743_o = setexecopc ? 1'b1 : n3742_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2098:82  */
  assign n3744_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2098:94  */
  assign n3746_o = n3744_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2098:73  */
  assign n3749_o = n3746_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3750_o = n3701_o ? make_berr : n3740_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3751_o = n3701_o & n3706_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3753_o = n3701_o ? n3718_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3755_o = n3701_o ? n3721_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3757_o = n3701_o ? n3724_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3759_o = n3701_o ? n3727_o : 1'b1;
  assign n3760_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3761_o = n3701_o ? n3760_o : n3743_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3763_o = n3701_o ? n3729_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3765_o = n3701_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2072:65  */
  assign n3766_o = n3701_o ? n3731_o : n3749_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3767_o = n3698_o ? n3750_o : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3768_o = n3698_o & n3751_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3770_o = n3698_o ? n3753_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3772_o = n3698_o ? n3755_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3774_o = n3698_o ? n3757_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3776_o = n3698_o ? n3759_o : 1'b0;
  assign n3777_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3778_o = n3698_o ? n3761_o : n3777_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3780_o = n3698_o ? n3763_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3782_o = n3698_o ? n3765_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2070:57  */
  assign n3784_o = n3698_o ? n3766_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2069:49  */
  assign n3786_o = n3568_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:66  */
  assign n3787_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:78  */
  assign n3789_o = n3787_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:74  */
  assign n3790_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:86  */
  assign n3792_o = n3790_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2109:75  */
  assign n3793_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2109:87  */
  assign n3795_o = n3793_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2109:105  */
  assign n3796_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2109:117  */
  assign n3798_o = n3796_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2109:96  */
  assign n3799_o = n3795_o | n3798_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:94  */
  assign n3800_o = n3792_o & n3799_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:101  */
  assign n3801_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:113  */
  assign n3803_o = n3801_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:91  */
  assign n3804_o = decodeopc & n3803_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:129  */
  assign n3806_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:148  */
  assign n3807_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:135  */
  assign n3808_o = n3806_o & n3807_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:120  */
  assign n3809_o = n3804_o | n3808_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2113:154  */
  assign n3810_o = n3809_o | direct_data;
  assign n3812_o = n1870_o[51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3813_o = n3883_o ? 1'b1 : n3812_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3815_o = n3875_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:65  */
  assign n3818_o = n3800_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:65  */
  assign n3821_o = n3800_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:65  */
  assign n3824_o = n3800_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:65  */
  assign n3827_o = n3800_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2108:65  */
  assign n3829_o = n3800_o & n3810_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:75  */
  assign n3830_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:87  */
  assign n3832_o = n3830_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2122:75  */
  assign n3833_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2122:87  */
  assign n3835_o = n3833_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2122:104  */
  assign n3836_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2122:116  */
  assign n3838_o = n3836_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2122:95  */
  assign n3839_o = n3835_o | n3838_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:95  */
  assign n3840_o = n3832_o & n3839_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2128:82  */
  assign n3843_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2128:94  */
  assign n3845_o = n3843_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2128:73  */
  assign n3848_o = n3845_o ? 1'b1 : 1'b0;
  assign n3850_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3851_o = n3868_o ? 1'b1 : n3850_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3854_o = n3840_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3857_o = n3840_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3860_o = n3840_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3863_o = n3840_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3866_o = n3840_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3868_o = n3840_o & setexecopc;
  assign n3869_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3870_o = n3840_o ? 1'b1 : n3869_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3872_o = n3840_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2121:65  */
  assign n3874_o = n3840_o ? n3848_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3875_o = n3789_o & n3800_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3877_o = n3789_o ? 1'b0 : n3854_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3878_o = n3789_o ? n3818_o : n3857_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3879_o = n3789_o ? n3821_o : n3860_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3880_o = n3789_o ? n3824_o : n3863_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3881_o = n3789_o ? n3827_o : n3866_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3883_o = n3789_o & n3829_o;
  assign n3884_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3885_o = n3789_o ? n3884_o : n3851_o;
  assign n3886_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3887_o = n3789_o ? n3886_o : n3870_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3889_o = n3789_o ? 1'b0 : n3872_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2107:57  */
  assign n3891_o = n3789_o ? 1'b0 : n3874_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2106:49  */
  assign n3893_o = n3568_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:66  */
  assign n3894_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:78  */
  assign n3896_o = n3894_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:74  */
  assign n3897_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:86  */
  assign n3899_o = n3897_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2142:75  */
  assign n3900_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2142:87  */
  assign n3902_o = n3900_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2142:105  */
  assign n3903_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2142:117  */
  assign n3905_o = n3903_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2142:96  */
  assign n3906_o = n3902_o | n3905_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:94  */
  assign n3907_o = n3899_o & n3906_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:109  */
  assign n3908_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:121  */
  assign n3910_o = n3908_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:99  */
  assign n3911_o = decodeopc & n3910_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:137  */
  assign n3913_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:156  */
  assign n3914_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:143  */
  assign n3915_o = n3913_o & n3914_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:128  */
  assign n3916_o = n3911_o | n3915_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2147:162  */
  assign n3917_o = n3916_o | direct_data;
  assign n3920_o = {1'b1, 1'b1};
  assign n3921_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n3922_o = n4023_o ? n3920_o : n3921_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:88  */
  assign n3923_o = exec[52];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:128  */
  assign n3924_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:140  */
  assign n3926_o = n3924_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:118  */
  assign n3927_o = decodeopc & n3926_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:100  */
  assign n3928_o = n3923_o | n3927_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:156  */
  assign n3930_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:175  */
  assign n3931_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:162  */
  assign n3932_o = n3930_o & n3931_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:147  */
  assign n3933_o = n3928_o | n3932_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2151:181  */
  assign n3934_o = n3933_o | direct_data;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n3936_o = n4012_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n3938_o = n4011_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2143:73  */
  assign n3939_o = svmode & n3934_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2143:73  */
  assign n3942_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2143:73  */
  assign n3945_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2143:73  */
  assign n3948_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2143:73  */
  assign n3951_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2143:73  */
  assign n3953_o = svmode & n3917_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3954_o = n3907_o & svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3955_o = n3907_o & n3939_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3957_o = n3907_o ? n3942_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3960_o = n3907_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3962_o = n3907_o ? n3945_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3964_o = n3907_o ? n3948_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3966_o = n3907_o ? n3951_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2141:65  */
  assign n3968_o = n3907_o & n3953_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:74  */
  assign n3969_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:86  */
  assign n3971_o = n3969_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2164:75  */
  assign n3972_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2164:87  */
  assign n3974_o = n3972_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2164:104  */
  assign n3975_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2164:116  */
  assign n3977_o = n3975_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2164:95  */
  assign n3978_o = n3974_o | n3977_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:94  */
  assign n3979_o = n3971_o & n3978_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2169:82  */
  assign n3982_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2169:94  */
  assign n3984_o = n3982_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2169:73  */
  assign n3987_o = n3984_o ? 1'b1 : 1'b0;
  assign n3989_o = n1870_o[53];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n3990_o = n4004_o ? 1'b1 : n3989_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n3993_o = n3979_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n3996_o = n3979_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n3999_o = n3979_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n4002_o = n3979_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n4004_o = n3979_o & setexecopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n4006_o = n3979_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n4008_o = n3979_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2163:65  */
  assign n4010_o = n3979_o ? n3987_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4011_o = n3896_o & n3954_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4012_o = n3896_o & n3955_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4014_o = n3896_o ? 1'b0 : n3993_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4016_o = n3896_o ? n3957_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4017_o = n3896_o ? n3960_o : n3996_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4019_o = n3896_o ? n3962_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4020_o = n3896_o ? n3964_o : n3999_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4021_o = n3896_o ? n3966_o : n4002_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4023_o = n3896_o & n3968_o;
  assign n4024_o = n1870_o[53];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4025_o = n3896_o ? n4024_o : n3990_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4027_o = n3896_o ? 1'b0 : n4006_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4029_o = n3896_o ? 1'b0 : n4008_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2140:57  */
  assign n4031_o = n3896_o ? 1'b0 : n4010_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2139:49  */
  assign n4033_o = n3568_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:66  */
  assign n4034_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:74  */
  assign n4035_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:86  */
  assign n4037_o = n4035_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:103  */
  assign n4038_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:107  */
  assign n4039_o = ~n4038_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:93  */
  assign n4040_o = n4037_o & n4039_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2187:82  */
  assign n4044_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2187:85  */
  assign n4045_o = ~n4044_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2187:73  */
  assign n4048_o = n4045_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2187:73  */
  assign n4050_o = n4045_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:83  */
  assign n4051_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:103  */
  assign n4052_o = opcode[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:120  */
  assign n4053_o = opcode[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:132  */
  assign n4055_o = n4053_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:111  */
  assign n4056_o = n4052_o | n4055_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2194:83  */
  assign n4057_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2194:95  */
  assign n4059_o = n4057_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2194:112  */
  assign n4060_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2194:124  */
  assign n4062_o = n4060_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2194:103  */
  assign n4063_o = n4059_o | n4062_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:139  */
  assign n4064_o = n4056_o & n4063_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:92  */
  assign n4065_o = n4051_o | n4064_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2195:83  */
  assign n4066_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2195:87  */
  assign n4067_o = ~n4066_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2195:102  */
  assign n4068_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2195:114  */
  assign n4070_o = n4068_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2196:82  */
  assign n4071_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2196:94  */
  assign n4073_o = n4071_o != 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2195:121  */
  assign n4074_o = n4070_o & n4073_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2197:82  */
  assign n4075_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2197:94  */
  assign n4077_o = n4075_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2196:102  */
  assign n4078_o = n4074_o & n4077_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2195:92  */
  assign n4079_o = n4067_o | n4078_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2194:133  */
  assign n4080_o = n4065_o & n4079_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2200:90  */
  assign n4082_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2200:93  */
  assign n4083_o = ~n4082_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4085_o = n4173_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:91  */
  assign n4086_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:103  */
  assign n4088_o = n4086_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:119  */
  assign n4089_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:131  */
  assign n4091_o = n4089_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:110  */
  assign n4092_o = n4088_o | n4091_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:148  */
  assign n4094_o = state == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:139  */
  assign n4095_o = n4092_o & n4094_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:81  */
  assign n4099_o = n4095_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2203:81  */
  assign n4101_o = n4095_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2207:90  */
  assign n4102_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2207:102  */
  assign n4104_o = n4102_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2207:81  */
  assign n4108_o = n4104_o ? 1'b1 : 1'b0;
  assign n4109_o = n1870_o[48];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2207:81  */
  assign n4110_o = n4104_o ? 1'b1 : n4109_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2211:89  */
  assign n4112_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2211:108  */
  assign n4113_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2211:95  */
  assign n4114_o = n4112_o & n4113_o;
  assign n4117_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4118_o = n4188_o ? 1'b1 : n4117_o;
  assign n4119_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4120_o = n4190_o ? 1'b1 : n4119_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:98  */
  assign n4122_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:110  */
  assign n4124_o = n4122_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:126  */
  assign n4125_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:138  */
  assign n4127_o = n4125_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:117  */
  assign n4128_o = n4124_o | n4127_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:154  */
  assign n4129_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:166  */
  assign n4131_o = n4129_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:145  */
  assign n4132_o = n4128_o | n4131_o;
  assign n4134_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:89  */
  assign n4135_o = n4132_o ? n4134_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2217:89  */
  assign n4138_o = n4132_o ? 7'b0011010 : 7'b0000001;
  assign n4139_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4140_o = n4194_o ? n4135_o : n4139_o;
  assign n4141_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4142_o = n4201_o ? 1'b1 : n4141_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2215:81  */
  assign n4143_o = decodeopc ? n4138_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2224:87  */
  assign n4144_o = set[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2227:106  */
  assign n4146_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2227:110  */
  assign n4147_o = ~n4146_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2227:97  */
  assign n4151_o = n4147_o ? 2'b11 : 2'b10;
  assign n4152_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4153_o = n4192_o ? 1'b1 : n4152_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2225:89  */
  assign n4156_o = movem_run ? n4151_o : 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2225:89  */
  assign n4158_o = movem_run & n4147_o;
  assign n4159_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4160_o = n4197_o ? 1'b1 : n4159_o;
  assign n4161_o = n1870_o[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4162_o = n4199_o ? 1'b1 : n4161_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2224:81  */
  assign n4164_o = n4172_o ? 7'b0011011 : n4143_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4165_o = n4174_o ? n4156_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2224:81  */
  assign n4167_o = n4144_o & n4158_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2224:81  */
  assign n4169_o = n4144_o & movem_run;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2224:81  */
  assign n4171_o = n4144_o & movem_run;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2224:81  */
  assign n4172_o = n4144_o & movem_run;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4173_o = n4080_o & n4083_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4174_o = n4080_o & n4144_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4177_o = n4080_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4179_o = n4080_o ? n4108_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4182_o = n4080_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4185_o = n4080_o ? 1'b0 : 1'b1;
  assign n4186_o = {1'b1, n4110_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4188_o = n4080_o & n4114_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4190_o = n4080_o & n4114_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4192_o = n4080_o & n4167_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4194_o = n4080_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4195_o = n4080_o ? n4186_o : n2136_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4197_o = n4080_o & n4169_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4199_o = n4080_o & n4171_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4201_o = n4080_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4203_o = n4080_o ? n4099_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4205_o = n4080_o ? n4101_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2193:73  */
  assign n4206_o = n4080_o ? n4164_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4207_o = n4040_o ? n4048_o : n4085_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4208_o = n4040_o ? n1985_o : n4165_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4210_o = n4040_o ? 1'b0 : n4177_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4213_o = n4040_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4215_o = n4040_o ? 1'b0 : n4179_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4217_o = n4040_o ? 1'b0 : n4182_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4219_o = n4040_o ? 1'b0 : n4185_o;
  assign n4220_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4221_o = n4040_o ? n4220_o : n4118_o;
  assign n4222_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4223_o = n4040_o ? n4222_o : n4120_o;
  assign n4224_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4225_o = n4040_o ? n4224_o : n4153_o;
  assign n4226_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4227_o = n4040_o ? n4226_o : n4140_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4228_o = n4040_o ? n2136_o : n4195_o;
  assign n4229_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4230_o = n4040_o ? n4229_o : n4160_o;
  assign n4231_o = n1870_o[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4232_o = n4040_o ? n4231_o : n4162_o;
  assign n4233_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4234_o = n4040_o ? n4233_o : n4142_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4236_o = n4040_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4238_o = n4040_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4240_o = n4040_o ? 1'b0 : n4203_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4241_o = n4040_o ? 1'b1 : n4205_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4243_o = n4040_o ? n4050_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2182:65  */
  assign n4244_o = n4040_o ? n2139_o : n4206_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:74  */
  assign n4245_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:82  */
  assign n4246_o = opcode[8:7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:94  */
  assign n4248_o = n4246_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:110  */
  assign n4249_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:122  */
  assign n4251_o = n4249_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:100  */
  assign n4252_o = n4248_o & n4251_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:141  */
  assign n4253_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:153  */
  assign n4255_o = n4253_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:171  */
  assign n4256_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:183  */
  assign n4258_o = n4256_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:162  */
  assign n4259_o = n4255_o | n4258_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:130  */
  assign n4260_o = n4252_o & n4259_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:190  */
  assign n4262_o = n4260_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2248:102  */
  assign n4263_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2248:105  */
  assign n4264_o = ~n4263_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2248:133  */
  assign n4265_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2248:141  */
  assign n4267_o = n4265_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2248:126  */
  assign n4269_o = 1'b0 | n4267_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2248:110  */
  assign n4270_o = n4264_o & n4269_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2248:91  */
  assign n4271_o = n4262_o & n4270_o;
  assign n4274_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2249:81  */
  assign n4275_o = decodeopc ? 1'b1 : n4274_o;
  assign n4276_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2249:81  */
  assign n4277_o = decodeopc ? 1'b1 : n4276_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2249:81  */
  assign n4279_o = decodeopc ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:96  */
  assign n4281_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:102  */
  assign n4282_o = n4281_o & nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:130  */
  assign n4283_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:142  */
  assign n4285_o = n4283_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:156  */
  assign n4286_o = exec[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:148  */
  assign n4287_o = n4285_o & n4286_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:120  */
  assign n4288_o = n4282_o | n4287_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2259:98  */
  assign n4291_o = sndopc[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:81  */
  assign n4293_o = n4299_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:81  */
  assign n4295_o = n4309_o ? 7'b1010100 : n4279_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:81  */
  assign n4299_o = n4288_o & n4291_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:81  */
  assign n4302_o = n4288_o ? 1'b1 : 1'b0;
  assign n4303_o = n1870_o[20];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4304_o = n4705_o ? 1'b1 : n4303_o;
  assign n4305_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4306_o = n4709_o ? 1'b1 : n4305_o;
  assign n4307_o = n1870_o[67];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4308_o = n4725_o ? 1'b1 : n4307_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2254:81  */
  assign n4309_o = n4288_o & n4291_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:85  */
  assign n4310_o = opcode[8:7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:97  */
  assign n4312_o = n4310_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:113  */
  assign n4313_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:125  */
  assign n4315_o = n4313_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:103  */
  assign n4316_o = n4312_o & n4315_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:144  */
  assign n4317_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:156  */
  assign n4319_o = n4317_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:174  */
  assign n4320_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:186  */
  assign n4322_o = n4320_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:165  */
  assign n4323_o = n4319_o | n4322_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:133  */
  assign n4324_o = n4316_o & n4323_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2270:84  */
  assign n4325_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2270:115  */
  assign n4326_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2270:123  */
  assign n4328_o = n4326_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2270:108  */
  assign n4330_o = 1'b0 | n4328_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2270:92  */
  assign n4331_o = n4325_o & n4330_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2271:83  */
  assign n4332_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2271:86  */
  assign n4333_o = ~n4332_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2271:114  */
  assign n4334_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2271:122  */
  assign n4336_o = n4334_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2271:107  */
  assign n4338_o = 1'b0 | n4336_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2271:91  */
  assign n4339_o = n4333_o & n4338_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2270:141  */
  assign n4340_o = n4331_o | n4339_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:193  */
  assign n4341_o = n4324_o & n4340_o;
  assign n4344_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4345_o = n4406_o ? 1'b1 : n4344_o;
  assign n4346_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4347_o = n4408_o ? 1'b1 : n4346_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2272:81  */
  assign n4349_o = decodeopc ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:96  */
  assign n4351_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:102  */
  assign n4352_o = n4351_o & nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:130  */
  assign n4353_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:142  */
  assign n4355_o = n4353_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:156  */
  assign n4356_o = exec[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:148  */
  assign n4357_o = n4355_o & n4356_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:120  */
  assign n4358_o = n4352_o | n4357_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2281:98  */
  assign n4359_o = opcode[6];
  assign n4361_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2281:89  */
  assign n4362_o = n4359_o ? n4361_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2281:89  */
  assign n4365_o = n4359_o ? 7'b1010101 : 7'b1010001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4367_o = n4387_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:81  */
  assign n4370_o = n4358_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:81  */
  assign n4373_o = n4358_o ? 1'b1 : 1'b0;
  assign n4374_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4375_o = n4404_o ? n4362_o : n4374_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2277:81  */
  assign n4376_o = n4358_o ? n4365_o : n4349_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2289:107  */
  assign n4377_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2289:119  */
  assign n4379_o = n4377_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2289:125  */
  assign n4380_o = n4379_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2289:97  */
  assign n4381_o = nextpass | n4380_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2289:81  */
  assign n4384_o = n4381_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4386_o = n4341_o ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4387_o = n4341_o & n4358_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4390_o = n4341_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4392_o = n4341_o ? n4370_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4394_o = n4341_o ? n4373_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4396_o = n4341_o ? n4384_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4399_o = n4341_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4402_o = n4341_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4404_o = n4341_o & n4358_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4406_o = n4341_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4408_o = n4341_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2269:73  */
  assign n4409_o = n4341_o ? n4376_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4411_o = n4271_o ? 2'b10 : n4386_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4412_o = n4271_o ? n4293_o : n4367_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4414_o = n4271_o ? 1'b1 : n4390_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4416_o = n4271_o ? 1'b0 : n4392_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4417_o = n4271_o ? n4302_o : n4394_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4419_o = n4271_o ? 1'b0 : n4396_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4421_o = n4271_o ? 1'b0 : n4399_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4423_o = n4271_o ? 1'b0 : n4402_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4425_o = n4271_o & n4288_o;
  assign n4426_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4427_o = n4271_o ? n4426_o : n4375_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4429_o = n4271_o & n4288_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4430_o = n4271_o ? n4275_o : n4345_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4432_o = n4271_o & n4288_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4433_o = n4271_o ? n4277_o : n4347_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2247:73  */
  assign n4434_o = n4271_o ? n4295_o : n4409_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:82  */
  assign n4435_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:90  */
  assign n4436_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:102  */
  assign n4438_o = n4436_o == 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:93  */
  assign n4441_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:105  */
  assign n4443_o = n4441_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:99  */
  assign n4444_o = opcode[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:116  */
  assign n4445_o = opcode[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:128  */
  assign n4447_o = n4445_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:107  */
  assign n4448_o = n4444_o | n4447_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2309:98  */
  assign n4449_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2309:110  */
  assign n4451_o = n4449_o != 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:135  */
  assign n4452_o = n4448_o & n4451_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2310:98  */
  assign n4453_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2310:110  */
  assign n4455_o = n4453_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2309:118  */
  assign n4456_o = n4452_o & n4455_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2313:128  */
  assign n4458_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2313:113  */
  assign n4459_o = nextpass & n4458_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2313:97  */
  assign n4462_o = n4459_o ? 2'b11 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4464_o = n4475_o ? 1'b1 : n1974_o;
  assign n4465_o = n2121_o[1];
  assign n4466_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4467_o = n1996_o ? n4465_o : n4466_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2313:97  */
  assign n4468_o = n4459_o ? 1'b1 : n4467_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4470_o = n4492_o ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2319:103  */
  assign n4471_o = set[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2319:97  */
  assign n4473_o = n4471_o ? 2'b01 : n4462_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4474_o = n4456_o ? n4473_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4475_o = n4456_o & n4459_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4478_o = n4456_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4481_o = n4456_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4484_o = n4456_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4487_o = n4456_o ? 1'b1 : 1'b0;
  assign n4488_o = n2121_o[1];
  assign n4489_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4490_o = n1996_o ? n4488_o : n4489_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4491_o = n4456_o ? n4468_o : n4490_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2308:89  */
  assign n4492_o = n4456_o & n4459_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4493_o = n4443_o ? n1985_o : n4474_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4494_o = n4443_o ? n1974_o : n4464_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4496_o = n4443_o ? 1'b0 : n4478_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4498_o = n4443_o ? 1'b1 : n4481_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4500_o = n4443_o ? 1'b1 : n4484_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4502_o = n4443_o ? 1'b0 : n4487_o;
  assign n4503_o = n2121_o[1];
  assign n4504_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4505_o = n1996_o ? n4503_o : n4504_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4506_o = n4443_o ? n4505_o : n4491_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2304:81  */
  assign n4507_o = n4443_o ? n2139_o : n4470_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4508_o = n4438_o ? n1985_o : n4493_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4509_o = n4438_o ? n1974_o : n4494_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4511_o = n4438_o ? 1'b0 : n4496_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4513_o = n4438_o ? 1'b0 : n4498_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4515_o = n4438_o ? 1'b0 : n4500_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4517_o = n4438_o ? 1'b0 : n4502_o;
  assign n4518_o = n2121_o[1];
  assign n4519_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4520_o = n1996_o ? n4518_o : n4519_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4521_o = n4438_o ? n4520_o : n4506_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4523_o = n4438_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4525_o = n4438_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2301:81  */
  assign n4526_o = n4438_o ? n2139_o : n4507_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:90  */
  assign n4527_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:102  */
  assign n4529_o = n4527_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4539_o = n4614_o ? 1'b1 : n1974_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2333:89  */
  assign n4542_o = decodeopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2333:89  */
  assign n4545_o = decodeopc ? 1'b1 : 1'b0;
  assign n4546_o = n1870_o[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4547_o = n4625_o ? 1'b1 : n4546_o;
  assign n4548_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4549_o = n4627_o ? 1'b1 : n4548_o;
  assign n4550_o = n2121_o[1];
  assign n4551_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4552_o = n1996_o ? n4550_o : n4551_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2333:89  */
  assign n4553_o = decodeopc ? 1'b1 : n4552_o;
  assign n4554_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4555_o = n4637_o ? 1'b1 : n4554_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4556_o = n4640_o ? 1'b1 : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4558_o = n4647_o ? 7'b0100011 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:98  */
  assign n4559_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:110  */
  assign n4561_o = n4559_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2346:99  */
  assign n4562_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2346:111  */
  assign n4564_o = n4562_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2346:128  */
  assign n4565_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2346:140  */
  assign n4567_o = n4565_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2346:119  */
  assign n4568_o = n4564_o | n4567_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:118  */
  assign n4569_o = n4561_o & n4568_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2354:106  */
  assign n4574_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2354:118  */
  assign n4576_o = n4574_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2354:97  */
  assign n4579_o = n4576_o ? 1'b1 : 1'b0;
  assign n4581_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4582_o = n4599_o ? 1'b1 : n4581_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4585_o = n4569_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4588_o = n4569_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4591_o = n4569_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4594_o = n4569_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4597_o = n4569_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4599_o = n4569_o & setexecopc;
  assign n4600_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4601_o = n4569_o ? 1'b1 : n4600_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4603_o = n4569_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4605_o = n4569_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4607_o = n4569_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2345:89  */
  assign n4609_o = n4569_o ? n4579_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4611_o = n4529_o ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4613_o = n4529_o ? 1'b0 : n4585_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4614_o = n4529_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4616_o = n4529_o ? n4542_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4617_o = n4529_o ? n4545_o : n4588_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4619_o = n4529_o ? 1'b0 : n4591_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4621_o = n4529_o ? 1'b0 : n4594_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4623_o = n4529_o ? 1'b0 : n4597_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4625_o = n4529_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4627_o = n4529_o & decodeopc;
  assign n4628_o = n2121_o[1];
  assign n4629_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4630_o = n1996_o ? n4628_o : n4629_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4631_o = n4529_o ? n4553_o : n4630_o;
  assign n4632_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4633_o = n4529_o ? 1'b1 : n4632_o;
  assign n4634_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4635_o = n4529_o ? n4634_o : n4582_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4637_o = n4529_o & decodeopc;
  assign n4638_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4639_o = n4529_o ? n4638_o : n4601_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4640_o = n4529_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4641_o = n4529_o ? 1'b1 : n4603_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4643_o = n4529_o ? 1'b0 : n4605_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4645_o = n4529_o ? 1'b0 : n4607_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4646_o = n4529_o ? 1'b1 : n4609_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2328:81  */
  assign n4647_o = n4529_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4649_o = n4435_o ? 2'b10 : n4611_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4650_o = n4435_o ? n4508_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4652_o = n4435_o ? 1'b0 : n4613_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4653_o = n4435_o ? n4509_o : n4539_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4655_o = n4435_o ? n4511_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4657_o = n4435_o ? 1'b0 : n4616_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4659_o = n4435_o ? 1'b0 : n4617_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4660_o = n4435_o ? n4513_o : n4619_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4661_o = n4435_o ? n4515_o : n4621_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4662_o = n4435_o ? n4517_o : n4623_o;
  assign n4663_o = {n4639_o, n4555_o, n4635_o};
  assign n4664_o = n1870_o[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4665_o = n4435_o ? n4664_o : n4547_o;
  assign n4666_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4667_o = n4435_o ? n4666_o : n4549_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4668_o = n4435_o ? n4521_o : n4631_o;
  assign n4669_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4670_o = n4435_o ? n4669_o : n4633_o;
  assign n4671_o = n1870_o[56:54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4672_o = n4435_o ? n4671_o : n4663_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4673_o = n4435_o ? n2130_o : n4556_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4675_o = n4435_o ? 1'b0 : n4641_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4677_o = n4435_o ? 1'b0 : n4643_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4679_o = n4435_o ? n4523_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4681_o = n4435_o ? 1'b0 : n4645_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4682_o = n4435_o ? n4525_o : n4646_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2299:73  */
  assign n4683_o = n4435_o ? n4526_o : n4558_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4684_o = n4245_o ? n4411_o : n4649_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4685_o = n4245_o ? n4412_o : n4650_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4687_o = n4245_o ? 1'b0 : n4652_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4688_o = n4245_o ? n1974_o : n4653_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4690_o = n4245_o ? 1'b0 : n4655_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4692_o = n4245_o ? 1'b0 : n4657_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4693_o = n4245_o ? n4414_o : n4659_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4695_o = n4245_o ? n4416_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4697_o = n4245_o ? n4417_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4699_o = n4245_o ? n4419_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4700_o = n4245_o ? n4421_o : n4660_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4701_o = n4245_o ? n4423_o : n4661_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4703_o = n4245_o ? 1'b0 : n4662_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4705_o = n4245_o & n4425_o;
  assign n4706_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4707_o = n4245_o ? n4427_o : n4706_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4709_o = n4245_o & n4429_o;
  assign n4710_o = n1870_o[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4711_o = n4245_o ? n4710_o : n4665_o;
  assign n4712_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4713_o = n4245_o ? n4430_o : n4712_o;
  assign n4714_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4715_o = n4245_o ? n4714_o : n4667_o;
  assign n4716_o = n2121_o[1];
  assign n4717_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4718_o = n1996_o ? n4716_o : n4717_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4719_o = n4245_o ? n4718_o : n4668_o;
  assign n4720_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4721_o = n4245_o ? n4720_o : n4670_o;
  assign n4722_o = n1870_o[56:54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4723_o = n4245_o ? n4722_o : n4672_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4725_o = n4245_o & n4432_o;
  assign n4726_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4727_o = n4245_o ? n4433_o : n4726_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4728_o = n4245_o ? n2130_o : n4673_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4730_o = n4245_o ? 1'b0 : n4675_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4732_o = n4245_o ? 1'b0 : n4677_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4734_o = n4245_o ? 1'b0 : n4679_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4736_o = n4245_o ? 1'b0 : n4681_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4738_o = n4245_o ? 1'b0 : n4682_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2245:65  */
  assign n4739_o = n4245_o ? n4434_o : n4683_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4740_o = n4034_o ? n4207_o : n4684_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4741_o = n4034_o ? n4208_o : n4685_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4743_o = n4034_o ? 1'b0 : n4687_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4744_o = n4034_o ? n1974_o : n4688_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4745_o = n4034_o ? n4210_o : n4690_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4747_o = n4034_o ? 1'b0 : n4692_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4748_o = n4034_o ? n4213_o : n4693_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4750_o = n4034_o ? 1'b0 : n4695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4752_o = n4034_o ? 1'b0 : n4697_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4754_o = n4034_o ? 1'b0 : n4699_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4756_o = n4034_o ? n4215_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4757_o = n4034_o ? n4217_o : n4700_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4758_o = n4034_o ? n4219_o : n4701_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4760_o = n4034_o ? 1'b0 : n4703_o;
  assign n4761_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4762_o = n4034_o ? n4221_o : n4761_o;
  assign n4763_o = n1870_o[20];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4764_o = n4034_o ? n4763_o : n4304_o;
  assign n4765_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4766_o = n4034_o ? n4765_o : n4707_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4767_o = n4034_o ? n4223_o : n4306_o;
  assign n4768_o = n1870_o[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4769_o = n4034_o ? n4768_o : n4711_o;
  assign n4770_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4771_o = n4034_o ? n4225_o : n4770_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4772_o = n4034_o ? n4227_o : n4713_o;
  assign n4773_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4774_o = n4034_o ? n4773_o : n4715_o;
  assign n4775_o = n2121_o[1];
  assign n4776_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4777_o = n1996_o ? n4775_o : n4776_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4778_o = n4034_o ? n4777_o : n4719_o;
  assign n4779_o = n4228_o[0];
  assign n4780_o = n1870_o[48];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4781_o = n4034_o ? n4779_o : n4780_o;
  assign n4782_o = n4228_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4783_o = n4034_o ? n4782_o : n4721_o;
  assign n4784_o = n4723_o[0];
  assign n4785_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4786_o = n4034_o ? n4785_o : n4784_o;
  assign n4787_o = n4723_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4788_o = n4034_o ? n4230_o : n4787_o;
  assign n4789_o = n4723_o[2];
  assign n4790_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4791_o = n4034_o ? n4790_o : n4789_o;
  assign n4792_o = n1870_o[67];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4793_o = n4034_o ? n4792_o : n4308_o;
  assign n4794_o = n1870_o[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4795_o = n4034_o ? n4232_o : n4794_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4796_o = n4034_o ? n4234_o : n4727_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4797_o = n4034_o ? n2130_o : n4728_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4799_o = n4034_o ? n4236_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4801_o = n4034_o ? 1'b0 : n4730_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4803_o = n4034_o ? n4238_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4805_o = n4034_o ? 1'b0 : n4732_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4807_o = n4034_o ? 1'b0 : n4734_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4809_o = n4034_o ? 1'b0 : n4736_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4811_o = n4034_o ? n4240_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4812_o = n4034_o ? n4241_o : n4738_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4814_o = n4034_o ? n4243_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2181:57  */
  assign n4815_o = n4034_o ? n4244_o : n4739_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2180:49  */
  assign n4817_o = n3568_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2180:59  */
  assign n4819_o = n3568_o == 3'b110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2180:59  */
  assign n4820_o = n4817_o | n4819_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:66  */
  assign n4821_o = opcode[7:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:78  */
  assign n4823_o = n4821_o == 5'b11111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:97  */
  assign n4824_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:109  */
  assign n4826_o = n4824_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:87  */
  assign n4827_o = n4823_o & n4826_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:75  */
  assign n4828_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:87  */
  assign n4830_o = n4828_o != 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2376:75  */
  assign n4831_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2376:87  */
  assign n4833_o = n4831_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2377:75  */
  assign n4834_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2377:87  */
  assign n4836_o = n4834_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2377:104  */
  assign n4837_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2377:116  */
  assign n4839_o = n4837_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2377:95  */
  assign n4840_o = n4836_o | n4839_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2376:95  */
  assign n4841_o = n4833_o & n4840_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:94  */
  assign n4842_o = n4830_o | n4841_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2378:76  */
  assign n4843_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2378:88  */
  assign n4845_o = n4843_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2378:105  */
  assign n4846_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2378:117  */
  assign n4848_o = n4846_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2378:95  */
  assign n4849_o = n4845_o | n4848_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2379:75  */
  assign n4850_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2379:87  */
  assign n4852_o = n4850_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2379:105  */
  assign n4853_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2379:117  */
  assign n4855_o = n4853_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2379:96  */
  assign n4856_o = n4852_o | n4855_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2378:127  */
  assign n4857_o = n4849_o & n4856_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2377:125  */
  assign n4858_o = n4842_o & n4857_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2383:90  */
  assign n4859_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2383:81  */
  assign n4862_o = n4859_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2381:73  */
  assign n4864_o = setexecopc ? n4862_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2381:73  */
  assign n4867_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2388:82  */
  assign n4869_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2388:94  */
  assign n4871_o = n4869_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2392:90  */
  assign n4872_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2392:102  */
  assign n4874_o = n4872_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2392:81  */
  assign n4877_o = n4874_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4879_o = n4888_o ? 2'b00 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2388:73  */
  assign n4882_o = n4871_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2388:73  */
  assign n4885_o = n4871_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2388:73  */
  assign n4887_o = n4871_o ? n4877_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4888_o = n4858_o & n4871_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4890_o = n4858_o ? n4882_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4892_o = n4858_o ? n4885_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4894_o = n4858_o ? n4864_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4896_o = n4858_o ? n4867_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4899_o = n4858_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4902_o = n4858_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4905_o = n4858_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4907_o = n4858_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2375:65  */
  assign n4909_o = n4858_o ? n4887_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4910_o = n4827_o ? n1882_o : n4879_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4912_o = n4827_o ? 1'b0 : n4890_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4914_o = n4827_o ? 1'b0 : n4892_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4916_o = n4827_o ? 1'b0 : n4894_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4918_o = n4827_o ? 1'b0 : n4896_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4920_o = n4827_o ? 1'b1 : n4899_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4922_o = n4827_o ? 1'b1 : n4902_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4924_o = n4827_o ? 1'b0 : n4905_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4926_o = n4827_o ? 1'b0 : n4907_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2371:57  */
  assign n4928_o = n4827_o ? 1'b0 : n4909_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2369:49  */
  assign n4930_o = n3568_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:66  */
  assign n4931_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:75  */
  assign n4932_o = opcode[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:92  */
  assign n4933_o = opcode[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:104  */
  assign n4935_o = n4933_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:83  */
  assign n4936_o = n4932_o | n4935_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2422:74  */
  assign n4937_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2422:86  */
  assign n4939_o = n4937_o != 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:111  */
  assign n4940_o = n4936_o & n4939_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2422:104  */
  assign n4941_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2422:116  */
  assign n4943_o = n4941_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2422:94  */
  assign n4944_o = n4940_o & n4943_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2426:80  */
  assign n4945_o = exec[63];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2426:73  */
  assign n4947_o = n4945_o ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:104  */
  assign n4949_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:89  */
  assign n4950_o = nextpass & n4949_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:120  */
  assign n4951_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:123  */
  assign n4952_o = ~n4951_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:110  */
  assign n4953_o = n4950_o & n4952_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:73  */
  assign n4956_o = n4953_o ? 2'b11 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n4958_o = n4994_o ? 1'b1 : n1974_o;
  assign n4959_o = n2121_o[1];
  assign n4960_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n4961_o = n1996_o ? n4959_o : n4960_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:73  */
  assign n4962_o = n4953_o ? 1'b1 : n4961_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2429:73  */
  assign n4964_o = n4953_o ? 7'b0011000 : n4947_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2436:87  */
  assign n4966_o = micro_state == 7'b0000101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2436:106  */
  assign n4967_o = brief[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2436:109  */
  assign n4968_o = ~n4967_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2436:97  */
  assign n4969_o = n4966_o & n4968_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2436:73  */
  assign n4971_o = n4969_o ? 1'b1 : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2439:81  */
  assign n4973_o = state == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2439:73  */
  assign n4976_o = n4973_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2443:79  */
  assign n4978_o = set[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2444:88  */
  assign n4979_o = exec[73];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2444:100  */
  assign n4980_o = ~n4979_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2444:105  */
  assign n4981_o = n4980_o | long_done;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2443:73  */
  assign n4983_o = n4985_o ? 1'b1 : n4971_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2443:73  */
  assign n4985_o = n4978_o & n4981_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2443:73  */
  assign n4987_o = n4978_o ? 2'b01 : n4956_o;
  assign n4988_o = n1870_o[63];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2443:73  */
  assign n4989_o = n4978_o ? 1'b1 : n4988_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n4990_o = n4944_o ? n4983_o : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n4992_o = n4944_o ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n4993_o = n4944_o ? n4987_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n4994_o = n4944_o & n4953_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n4996_o = n4944_o ? n4976_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n4999_o = n4944_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n5002_o = n4944_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n5005_o = n4944_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n5008_o = n4944_o ? 1'b1 : 1'b0;
  assign n5009_o = {1'b1, n4989_o};
  assign n5010_o = n2121_o[1];
  assign n5011_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5012_o = n1996_o ? n5010_o : n5011_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n5013_o = n4944_o ? n4962_o : n5012_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5014_o = n5562_o ? n5009_o : n2137_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2421:65  */
  assign n5015_o = n4944_o ? n4964_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:76  */
  assign n5016_o = opcode[6:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:73  */
  assign n5018_o = n5016_o == 7'b1000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:87  */
  assign n5020_o = n5016_o == 7'b1000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:87  */
  assign n5021_o = n5018_o | n5020_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:97  */
  assign n5023_o = n5016_o == 7'b1000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:97  */
  assign n5024_o = n5021_o | n5023_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:107  */
  assign n5026_o = n5016_o == 7'b1000011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:107  */
  assign n5027_o = n5024_o | n5026_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:117  */
  assign n5029_o = n5016_o == 7'b1000100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:117  */
  assign n5030_o = n5027_o | n5029_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:127  */
  assign n5032_o = n5016_o == 7'b1000101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:127  */
  assign n5033_o = n5030_o | n5032_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:137  */
  assign n5035_o = n5016_o == 7'b1000110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:137  */
  assign n5036_o = n5033_o | n5035_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:147  */
  assign n5038_o = n5016_o == 7'b1000111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:147  */
  assign n5039_o = n5036_o | n5038_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:157  */
  assign n5041_o = n5016_o == 7'b1001000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2456:157  */
  assign n5042_o = n5039_o | n5041_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:87  */
  assign n5044_o = n5016_o == 7'b1001001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:87  */
  assign n5045_o = n5042_o | n5044_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:97  */
  assign n5047_o = n5016_o == 7'b1001010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:97  */
  assign n5048_o = n5045_o | n5047_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:107  */
  assign n5050_o = n5016_o == 7'b1001011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:107  */
  assign n5051_o = n5048_o | n5050_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:117  */
  assign n5053_o = n5016_o == 7'b1001100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:117  */
  assign n5054_o = n5051_o | n5053_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:127  */
  assign n5056_o = n5016_o == 7'b1001101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:127  */
  assign n5057_o = n5054_o | n5056_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:137  */
  assign n5059_o = n5016_o == 7'b1001110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:137  */
  assign n5060_o = n5057_o | n5059_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:147  */
  assign n5062_o = n5016_o == 7'b1001111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2457:147  */
  assign n5063_o = n5060_o | n5062_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2466:81  */
  assign n5071_o = decodeopc ? 1'b1 : n1974_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2466:81  */
  assign n5074_o = decodeopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2466:81  */
  assign n5077_o = decodeopc ? 1'b1 : 1'b0;
  assign n5078_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2466:81  */
  assign n5079_o = decodeopc ? 1'b1 : n5078_o;
  assign n5080_o = n2121_o[1];
  assign n5081_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5082_o = n1996_o ? n5080_o : n5081_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2466:81  */
  assign n5083_o = decodeopc ? 1'b1 : n5082_o;
  assign n5084_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2466:81  */
  assign n5085_o = decodeopc ? 1'b1 : n5084_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2466:81  */
  assign n5087_o = decodeopc ? 7'b0100011 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:73  */
  assign n5089_o = n5016_o == 7'b1010000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:87  */
  assign n5091_o = n5016_o == 7'b1010001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:87  */
  assign n5092_o = n5089_o | n5091_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:97  */
  assign n5094_o = n5016_o == 7'b1010010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:97  */
  assign n5095_o = n5092_o | n5094_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:107  */
  assign n5097_o = n5016_o == 7'b1010011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:107  */
  assign n5098_o = n5095_o | n5097_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:117  */
  assign n5100_o = n5016_o == 7'b1010100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:117  */
  assign n5101_o = n5098_o | n5100_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:127  */
  assign n5103_o = n5016_o == 7'b1010101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:127  */
  assign n5104_o = n5101_o | n5103_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:137  */
  assign n5106_o = n5016_o == 7'b1010110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:137  */
  assign n5107_o = n5104_o | n5106_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:147  */
  assign n5109_o = n5016_o == 7'b1010111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2461:147  */
  assign n5110_o = n5107_o | n5109_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2481:81  */
  assign n5117_o = decodeopc ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2481:81  */
  assign n5119_o = decodeopc ? 1'b1 : n1974_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2481:81  */
  assign n5122_o = decodeopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2481:81  */
  assign n5125_o = decodeopc ? 1'b1 : 1'b0;
  assign n5126_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2481:81  */
  assign n5127_o = decodeopc ? 1'b1 : n5126_o;
  assign n5128_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2481:81  */
  assign n5129_o = decodeopc ? 1'b1 : n5128_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2481:81  */
  assign n5131_o = decodeopc ? 7'b0100101 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:73  */
  assign n5133_o = n5016_o == 7'b1011000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:87  */
  assign n5135_o = n5016_o == 7'b1011001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:87  */
  assign n5136_o = n5133_o | n5135_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:97  */
  assign n5138_o = n5016_o == 7'b1011010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:97  */
  assign n5139_o = n5136_o | n5138_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:107  */
  assign n5141_o = n5016_o == 7'b1011011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:107  */
  assign n5142_o = n5139_o | n5141_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:117  */
  assign n5144_o = n5016_o == 7'b1011100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:117  */
  assign n5145_o = n5142_o | n5144_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:127  */
  assign n5147_o = n5016_o == 7'b1011101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:127  */
  assign n5148_o = n5145_o | n5147_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:137  */
  assign n5150_o = n5016_o == 7'b1011110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:137  */
  assign n5151_o = n5148_o | n5150_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:147  */
  assign n5153_o = n5016_o == 7'b1011111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2476:147  */
  assign n5154_o = n5151_o | n5153_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2492:81  */
  assign n5157_o = svmode ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2492:81  */
  assign n5160_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2492:81  */
  assign n5163_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2492:81  */
  assign n5166_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2492:81  */
  assign n5169_o = svmode ? 1'b0 : 1'b1;
  assign n5170_o = n1976_o[0];
  assign n5171_o = n1870_o[65];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:17  */
  assign n5172_o = n1969_o ? n5170_o : n5171_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2492:81  */
  assign n5173_o = svmode ? 1'b1 : n5172_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:73  */
  assign n5175_o = n5016_o == 7'b1100000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:87  */
  assign n5177_o = n5016_o == 7'b1100001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:87  */
  assign n5178_o = n5175_o | n5177_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:97  */
  assign n5180_o = n5016_o == 7'b1100010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:97  */
  assign n5181_o = n5178_o | n5180_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:107  */
  assign n5183_o = n5016_o == 7'b1100011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:107  */
  assign n5184_o = n5181_o | n5183_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:117  */
  assign n5186_o = n5016_o == 7'b1100100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:117  */
  assign n5187_o = n5184_o | n5186_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:127  */
  assign n5189_o = n5016_o == 7'b1100101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:127  */
  assign n5190_o = n5187_o | n5189_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:137  */
  assign n5192_o = n5016_o == 7'b1100110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:137  */
  assign n5193_o = n5190_o | n5192_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:147  */
  assign n5195_o = n5016_o == 7'b1100111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2491:147  */
  assign n5196_o = n5193_o | n5195_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2504:81  */
  assign n5200_o = svmode ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2504:81  */
  assign n5203_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2504:81  */
  assign n5206_o = svmode ? 1'b0 : 1'b1;
  assign n5207_o = n1976_o[1];
  assign n5208_o = n1870_o[66];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:17  */
  assign n5209_o = n1969_o ? n5207_o : n5208_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2504:81  */
  assign n5210_o = svmode ? 1'b1 : n5209_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2504:81  */
  assign n5212_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:73  */
  assign n5214_o = n5016_o == 7'b1101000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:87  */
  assign n5216_o = n5016_o == 7'b1101001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:87  */
  assign n5217_o = n5214_o | n5216_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:97  */
  assign n5219_o = n5016_o == 7'b1101010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:97  */
  assign n5220_o = n5217_o | n5219_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:107  */
  assign n5222_o = n5016_o == 7'b1101011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:107  */
  assign n5223_o = n5220_o | n5222_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:117  */
  assign n5225_o = n5016_o == 7'b1101100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:117  */
  assign n5226_o = n5223_o | n5225_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:127  */
  assign n5228_o = n5016_o == 7'b1101101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:127  */
  assign n5229_o = n5226_o | n5228_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:137  */
  assign n5231_o = n5016_o == 7'b1101110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:137  */
  assign n5232_o = n5229_o | n5231_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:147  */
  assign n5234_o = n5016_o == 7'b1101111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2503:147  */
  assign n5235_o = n5232_o | n5234_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2515:90  */
  assign n5236_o = ~svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2520:89  */
  assign n5240_o = decodeopc ? 6'b000000 : n1867_o;
  assign n5241_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2520:89  */
  assign n5242_o = decodeopc ? 1'b1 : n5241_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2515:81  */
  assign n5243_o = n5236_o ? n1867_o : n5240_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2515:81  */
  assign n5246_o = n5236_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2515:81  */
  assign n5249_o = n5236_o ? 1'b1 : 1'b0;
  assign n5250_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2515:81  */
  assign n5251_o = n5236_o ? n5250_o : n5242_o;
  assign n5252_o = n1870_o[74];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2515:81  */
  assign n5253_o = n5236_o ? n5252_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2514:73  */
  assign n5255_o = n5016_o == 7'b1110000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2526:73  */
  assign n5257_o = n5016_o == 7'b1110001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2529:90  */
  assign n5258_o = ~svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2533:89  */
  assign n5260_o = decodeopc ? 1'b1 : n2107_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2533:89  */
  assign n5263_o = decodeopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2537:89  */
  assign n5265_o = stop ? 1'b1 : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2529:81  */
  assign n5266_o = n5258_o ? make_berr : n5265_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2529:81  */
  assign n5267_o = n5258_o ? n2107_o : n5260_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2529:81  */
  assign n5270_o = n5258_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2529:81  */
  assign n5273_o = n5258_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2529:81  */
  assign n5275_o = n5258_o ? 1'b0 : n5263_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2528:73  */
  assign n5277_o = n5016_o == 7'b1110010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:104  */
  assign n5278_o = opcode[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:95  */
  assign n5279_o = svmode | n5278_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2549:106  */
  assign n5281_o = opcode[2];
  assign n5284_o = n1870_o[59];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2549:97  */
  assign n5285_o = n5281_o ? n5284_o : 1'b1;
  assign n5286_o = n1870_o[60];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2549:97  */
  assign n5287_o = n5281_o ? 1'b1 : n5286_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5289_o = n5301_o ? 2'b10 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5291_o = n5302_o ? 1'b1 : n1974_o;
  assign n5292_o = {n5287_o, n5285_o};
  assign n5293_o = n2121_o[0];
  assign n5294_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5295_o = n1996_o ? n5293_o : n5294_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2545:89  */
  assign n5296_o = decodeopc ? 1'b1 : n5295_o;
  assign n5297_o = n1870_o[60:59];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5298_o = n5314_o ? n5292_o : n5297_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5300_o = n5315_o ? 7'b0101011 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5301_o = n5279_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5302_o = n5279_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5305_o = n5279_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5308_o = n5279_o ? 1'b0 : 1'b1;
  assign n5309_o = n2121_o[0];
  assign n5310_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5311_o = n1996_o ? n5309_o : n5310_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5312_o = n5279_o ? n5296_o : n5311_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5314_o = n5279_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2544:81  */
  assign n5315_o = n5279_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2543:73  */
  assign n5317_o = n5016_o == 7'b1110011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2543:87  */
  assign n5319_o = n5016_o == 7'b1110111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2543:87  */
  assign n5320_o = n5317_o | n5319_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2563:81  */
  assign n5325_o = decodeopc ? 2'b10 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2563:81  */
  assign n5327_o = decodeopc ? 1'b1 : n1974_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2563:81  */
  assign n5329_o = decodeopc ? 1'b1 : n2113_o;
  assign n5330_o = {1'b1, 1'b1};
  assign n5331_o = n2121_o[0];
  assign n5332_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5333_o = n1996_o ? n5331_o : n5332_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2563:81  */
  assign n5334_o = decodeopc ? 1'b1 : n5333_o;
  assign n5335_o = n1870_o[58:57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2563:81  */
  assign n5336_o = decodeopc ? n5330_o : n5335_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2563:81  */
  assign n5338_o = decodeopc ? 7'b0110000 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2561:73  */
  assign n5340_o = n5016_o == 7'b1110100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2576:81  */
  assign n5345_o = decodeopc ? 2'b10 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2576:81  */
  assign n5347_o = decodeopc ? 1'b1 : n1974_o;
  assign n5348_o = {1'b1, 1'b1};
  assign n5349_o = n2121_o[0];
  assign n5350_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5351_o = n1996_o ? n5349_o : n5350_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2576:81  */
  assign n5352_o = decodeopc ? 1'b1 : n5351_o;
  assign n5353_o = n1870_o[58:57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2576:81  */
  assign n5354_o = decodeopc ? n5348_o : n5353_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2576:81  */
  assign n5356_o = decodeopc ? 7'b0011000 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2574:73  */
  assign n5358_o = n5016_o == 7'b1110101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2586:81  */
  assign n5360_o = decodeopc ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2589:89  */
  assign n5361_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2589:106  */
  assign n5363_o = state == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2589:97  */
  assign n5364_o = n5361_o & n5363_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2589:81  */
  assign n5367_o = n5364_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2589:81  */
  assign n5370_o = n5364_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2585:73  */
  assign n5372_o = n5016_o == 7'b1110110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:87  */
  assign n5374_o = cpu == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:93  */
  assign n5375_o = ~svmode;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2603:106  */
  assign n5376_o = last_data_read[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2603:119  */
  assign n5378_o = n5376_o == 12'b100000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2605:106  */
  assign n5380_o = opcode[0];
  assign n5382_o = n1976_o[0];
  assign n5383_o = n1870_o[65];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:17  */
  assign n5384_o = n1969_o ? n5382_o : n5383_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2605:97  */
  assign n5385_o = n5380_o ? 1'b1 : n5384_o;
  assign n5386_o = {1'b1, n5385_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2603:89  */
  assign n5387_o = n5378_o ? n5386_o : n1978_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2609:98  */
  assign n5388_o = opcode[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2609:101  */
  assign n5389_o = ~n5388_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2609:89  */
  assign n5393_o = n5389_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2609:89  */
  assign n5395_o = n5389_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2614:89  */
  assign n5397_o = decodeopc ? 1'b1 : n2110_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2614:89  */
  assign n5399_o = decodeopc ? 7'b1001001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:81  */
  assign n5401_o = n5375_o ? n1882_o : 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:81  */
  assign n5402_o = n5375_o ? n2110_o : n5397_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:81  */
  assign n5405_o = n5375_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:81  */
  assign n5408_o = n5375_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:81  */
  assign n5409_o = n5375_o ? n1978_o : n5387_o;
  assign n5410_o = {n5395_o, n5393_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:81  */
  assign n5412_o = n5375_o ? 2'b00 : n5410_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2598:81  */
  assign n5413_o = n5375_o ? n2139_o : n5399_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5414_o = n5374_o ? n1882_o : n5401_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5415_o = n5374_o ? n2110_o : n5402_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5418_o = n5374_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5420_o = n5374_o ? 1'b0 : n5405_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5422_o = n5374_o ? 1'b1 : n5408_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5423_o = n5374_o ? n1978_o : n5409_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5425_o = n5374_o ? 2'b00 : n5412_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2595:81  */
  assign n5426_o = n5374_o ? n2139_o : n5413_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2594:73  */
  assign n5428_o = n5016_o == 7'b1111010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2594:87  */
  assign n5430_o = n5016_o == 7'b1111011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2594:87  */
  assign n5431_o = n5428_o | n5430_o;
  assign n5432_o = {n5431_o, n5372_o, n5358_o, n5340_o, n5320_o, n5277_o, n5257_o, n5255_o, n5235_o, n5196_o, n5154_o, n5110_o, n5063_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5433_o = make_berr;
      13'b0100000000000: n5433_o = make_berr;
      13'b0010000000000: n5433_o = make_berr;
      13'b0001000000000: n5433_o = make_berr;
      13'b0000100000000: n5433_o = make_berr;
      13'b0000010000000: n5433_o = n5266_o;
      13'b0000001000000: n5433_o = make_berr;
      13'b0000000100000: n5433_o = make_berr;
      13'b0000000010000: n5433_o = make_berr;
      13'b0000000001000: n5433_o = make_berr;
      13'b0000000000100: n5433_o = make_berr;
      13'b0000000000010: n5433_o = make_berr;
      13'b0000000000001: n5433_o = make_berr;
      default: n5433_o = make_berr;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5438_o = n5414_o;
      13'b0100000000000: n5438_o = n1882_o;
      13'b0010000000000: n5438_o = 2'b10;
      13'b0001000000000: n5438_o = 2'b10;
      13'b0000100000000: n5438_o = n1882_o;
      13'b0000010000000: n5438_o = n1882_o;
      13'b0000001000000: n5438_o = n1882_o;
      13'b0000000100000: n5438_o = n1882_o;
      13'b0000000010000: n5438_o = n5200_o;
      13'b0000000001000: n5438_o = n5157_o;
      13'b0000000000100: n5438_o = 2'b10;
      13'b0000000000010: n5438_o = 2'b10;
      13'b0000000000001: n5438_o = n1882_o;
      default: n5438_o = n1882_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5439_o = n1985_o;
      13'b0100000000000: n5439_o = n5360_o;
      13'b0010000000000: n5439_o = n5345_o;
      13'b0001000000000: n5439_o = n5325_o;
      13'b0000100000000: n5439_o = n5289_o;
      13'b0000010000000: n5439_o = n1985_o;
      13'b0000001000000: n5439_o = n1985_o;
      13'b0000000100000: n5439_o = n1985_o;
      13'b0000000010000: n5439_o = n1985_o;
      13'b0000000001000: n5439_o = n1985_o;
      13'b0000000000100: n5439_o = n5117_o;
      13'b0000000000010: n5439_o = n1985_o;
      13'b0000000000001: n5439_o = n1985_o;
      default: n5439_o = n1985_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5440_o = n2107_o;
      13'b0100000000000: n5440_o = n2107_o;
      13'b0010000000000: n5440_o = n2107_o;
      13'b0001000000000: n5440_o = n2107_o;
      13'b0000100000000: n5440_o = n2107_o;
      13'b0000010000000: n5440_o = n5267_o;
      13'b0000001000000: n5440_o = n2107_o;
      13'b0000000100000: n5440_o = n2107_o;
      13'b0000000010000: n5440_o = n2107_o;
      13'b0000000001000: n5440_o = n2107_o;
      13'b0000000000100: n5440_o = n2107_o;
      13'b0000000000010: n5440_o = n2107_o;
      13'b0000000000001: n5440_o = n2107_o;
      default: n5440_o = n2107_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5441_o = n5415_o;
      13'b0100000000000: n5441_o = n2110_o;
      13'b0010000000000: n5441_o = n2110_o;
      13'b0001000000000: n5441_o = n2110_o;
      13'b0000100000000: n5441_o = n2110_o;
      13'b0000010000000: n5441_o = n2110_o;
      13'b0000001000000: n5441_o = n2110_o;
      13'b0000000100000: n5441_o = n2110_o;
      13'b0000000010000: n5441_o = n2110_o;
      13'b0000000001000: n5441_o = n2110_o;
      13'b0000000000100: n5441_o = n2110_o;
      13'b0000000000010: n5441_o = n2110_o;
      13'b0000000000001: n5441_o = n2110_o;
      default: n5441_o = n2110_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5442_o = n1974_o;
      13'b0100000000000: n5442_o = n1974_o;
      13'b0010000000000: n5442_o = n5347_o;
      13'b0001000000000: n5442_o = n5327_o;
      13'b0000100000000: n5442_o = n5291_o;
      13'b0000010000000: n5442_o = n1974_o;
      13'b0000001000000: n5442_o = n1974_o;
      13'b0000000100000: n5442_o = n1974_o;
      13'b0000000010000: n5442_o = n1974_o;
      13'b0000000001000: n5442_o = n1974_o;
      13'b0000000000100: n5442_o = n5119_o;
      13'b0000000000010: n5442_o = n5071_o;
      13'b0000000000001: n5442_o = n1974_o;
      default: n5442_o = n1974_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5444_o = 1'b0;
      13'b0100000000000: n5444_o = 1'b0;
      13'b0010000000000: n5444_o = 1'b0;
      13'b0001000000000: n5444_o = 1'b0;
      13'b0000100000000: n5444_o = 1'b0;
      13'b0000010000000: n5444_o = 1'b0;
      13'b0000001000000: n5444_o = 1'b0;
      13'b0000000100000: n5444_o = 1'b0;
      13'b0000000010000: n5444_o = 1'b0;
      13'b0000000001000: n5444_o = n5160_o;
      13'b0000000000100: n5444_o = n5122_o;
      13'b0000000000010: n5444_o = n5074_o;
      13'b0000000000001: n5444_o = 1'b0;
      default: n5444_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5446_o = 1'b0;
      13'b0100000000000: n5446_o = 1'b0;
      13'b0010000000000: n5446_o = 1'b0;
      13'b0001000000000: n5446_o = 1'b0;
      13'b0000100000000: n5446_o = 1'b0;
      13'b0000010000000: n5446_o = 1'b0;
      13'b0000001000000: n5446_o = 1'b0;
      13'b0000000100000: n5446_o = 1'b0;
      13'b0000000010000: n5446_o = 1'b0;
      13'b0000000001000: n5446_o = n5163_o;
      13'b0000000000100: n5446_o = n5125_o;
      13'b0000000000010: n5446_o = n5077_o;
      13'b0000000000001: n5446_o = 1'b0;
      default: n5446_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5447_o = n1867_o;
      13'b0100000000000: n5447_o = n1867_o;
      13'b0010000000000: n5447_o = n1867_o;
      13'b0001000000000: n5447_o = n1867_o;
      13'b0000100000000: n5447_o = n1867_o;
      13'b0000010000000: n5447_o = n1867_o;
      13'b0000001000000: n5447_o = n1867_o;
      13'b0000000100000: n5447_o = n5243_o;
      13'b0000000010000: n5447_o = n1867_o;
      13'b0000000001000: n5447_o = n1867_o;
      13'b0000000000100: n5447_o = n1867_o;
      13'b0000000000010: n5447_o = n1867_o;
      13'b0000000000001: n5447_o = n1867_o;
      default: n5447_o = n1867_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5448_o = n2113_o;
      13'b0100000000000: n5448_o = n2113_o;
      13'b0010000000000: n5448_o = n2113_o;
      13'b0001000000000: n5448_o = n5329_o;
      13'b0000100000000: n5448_o = n2113_o;
      13'b0000010000000: n5448_o = n2113_o;
      13'b0000001000000: n5448_o = n2113_o;
      13'b0000000100000: n5448_o = n2113_o;
      13'b0000000010000: n5448_o = n2113_o;
      13'b0000000001000: n5448_o = n2113_o;
      13'b0000000000100: n5448_o = n2113_o;
      13'b0000000000010: n5448_o = n2113_o;
      13'b0000000000001: n5448_o = n2113_o;
      default: n5448_o = n2113_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5451_o = n5418_o;
      13'b0100000000000: n5451_o = 1'b0;
      13'b0010000000000: n5451_o = 1'b0;
      13'b0001000000000: n5451_o = 1'b0;
      13'b0000100000000: n5451_o = 1'b0;
      13'b0000010000000: n5451_o = 1'b0;
      13'b0000001000000: n5451_o = 1'b0;
      13'b0000000100000: n5451_o = 1'b0;
      13'b0000000010000: n5451_o = 1'b0;
      13'b0000000001000: n5451_o = 1'b0;
      13'b0000000000100: n5451_o = 1'b0;
      13'b0000000000010: n5451_o = 1'b0;
      13'b0000000000001: n5451_o = 1'b0;
      default: n5451_o = 1'b1;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5453_o = n5420_o;
      13'b0100000000000: n5453_o = 1'b0;
      13'b0010000000000: n5453_o = 1'b0;
      13'b0001000000000: n5453_o = 1'b0;
      13'b0000100000000: n5453_o = n5305_o;
      13'b0000010000000: n5453_o = n5270_o;
      13'b0000001000000: n5453_o = 1'b0;
      13'b0000000100000: n5453_o = n5246_o;
      13'b0000000010000: n5453_o = n5203_o;
      13'b0000000001000: n5453_o = n5166_o;
      13'b0000000000100: n5453_o = 1'b0;
      13'b0000000000010: n5453_o = 1'b0;
      13'b0000000000001: n5453_o = 1'b0;
      default: n5453_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5456_o = 1'b0;
      13'b0100000000000: n5456_o = 1'b0;
      13'b0010000000000: n5456_o = 1'b0;
      13'b0001000000000: n5456_o = 1'b0;
      13'b0000100000000: n5456_o = 1'b0;
      13'b0000010000000: n5456_o = 1'b0;
      13'b0000001000000: n5456_o = 1'b0;
      13'b0000000100000: n5456_o = 1'b0;
      13'b0000000010000: n5456_o = 1'b0;
      13'b0000000001000: n5456_o = 1'b0;
      13'b0000000000100: n5456_o = 1'b0;
      13'b0000000000010: n5456_o = 1'b0;
      13'b0000000000001: n5456_o = 1'b1;
      default: n5456_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5458_o = 1'b0;
      13'b0100000000000: n5458_o = n5367_o;
      13'b0010000000000: n5458_o = 1'b0;
      13'b0001000000000: n5458_o = 1'b0;
      13'b0000100000000: n5458_o = 1'b0;
      13'b0000010000000: n5458_o = 1'b0;
      13'b0000001000000: n5458_o = 1'b0;
      13'b0000000100000: n5458_o = 1'b0;
      13'b0000000010000: n5458_o = 1'b0;
      13'b0000000001000: n5458_o = 1'b0;
      13'b0000000000100: n5458_o = 1'b0;
      13'b0000000000010: n5458_o = 1'b0;
      13'b0000000000001: n5458_o = 1'b0;
      default: n5458_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5462_o = n5422_o;
      13'b0100000000000: n5462_o = n5370_o;
      13'b0010000000000: n5462_o = 1'b0;
      13'b0001000000000: n5462_o = 1'b0;
      13'b0000100000000: n5462_o = n5308_o;
      13'b0000010000000: n5462_o = n5273_o;
      13'b0000001000000: n5462_o = 1'b0;
      13'b0000000100000: n5462_o = n5249_o;
      13'b0000000010000: n5462_o = n5206_o;
      13'b0000000001000: n5462_o = n5169_o;
      13'b0000000000100: n5462_o = 1'b0;
      13'b0000000000010: n5462_o = 1'b0;
      13'b0000000000001: n5462_o = 1'b1;
      default: n5462_o = 1'b1;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5464_o = 1'b0;
      13'b0100000000000: n5464_o = 1'b0;
      13'b0010000000000: n5464_o = 1'b0;
      13'b0001000000000: n5464_o = 1'b0;
      13'b0000100000000: n5464_o = 1'b0;
      13'b0000010000000: n5464_o = n5275_o;
      13'b0000001000000: n5464_o = 1'b0;
      13'b0000000100000: n5464_o = 1'b0;
      13'b0000000010000: n5464_o = 1'b0;
      13'b0000000001000: n5464_o = 1'b0;
      13'b0000000000100: n5464_o = 1'b0;
      13'b0000000000010: n5464_o = 1'b0;
      13'b0000000000001: n5464_o = 1'b0;
      default: n5464_o = 1'b0;
    endcase
  assign n5465_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5466_o = n5465_o;
      13'b0100000000000: n5466_o = n5465_o;
      13'b0010000000000: n5466_o = n5465_o;
      13'b0001000000000: n5466_o = n5465_o;
      13'b0000100000000: n5466_o = n5465_o;
      13'b0000010000000: n5466_o = n5465_o;
      13'b0000001000000: n5466_o = n5465_o;
      13'b0000000100000: n5466_o = n5465_o;
      13'b0000000010000: n5466_o = n5465_o;
      13'b0000000001000: n5466_o = n5465_o;
      13'b0000000000100: n5466_o = n5127_o;
      13'b0000000000010: n5466_o = n5465_o;
      13'b0000000000001: n5466_o = n5465_o;
      default: n5466_o = n5465_o;
    endcase
  assign n5467_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5468_o = n5467_o;
      13'b0100000000000: n5468_o = n5467_o;
      13'b0010000000000: n5468_o = n5467_o;
      13'b0001000000000: n5468_o = n5467_o;
      13'b0000100000000: n5468_o = n5467_o;
      13'b0000010000000: n5468_o = n5467_o;
      13'b0000001000000: n5468_o = n5467_o;
      13'b0000000100000: n5468_o = n5251_o;
      13'b0000000010000: n5468_o = n5467_o;
      13'b0000000001000: n5468_o = n5467_o;
      13'b0000000000100: n5468_o = n5467_o;
      13'b0000000000010: n5468_o = n5467_o;
      13'b0000000000001: n5468_o = n5467_o;
      default: n5468_o = n5467_o;
    endcase
  assign n5469_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5470_o = n5469_o;
      13'b0100000000000: n5470_o = n5469_o;
      13'b0010000000000: n5470_o = n5469_o;
      13'b0001000000000: n5470_o = n5469_o;
      13'b0000100000000: n5470_o = n5469_o;
      13'b0000010000000: n5470_o = n5469_o;
      13'b0000001000000: n5470_o = n5469_o;
      13'b0000000100000: n5470_o = n5469_o;
      13'b0000000010000: n5470_o = n5469_o;
      13'b0000000001000: n5470_o = n5469_o;
      13'b0000000000100: n5470_o = n5129_o;
      13'b0000000000010: n5470_o = n5469_o;
      13'b0000000000001: n5470_o = n5469_o;
      default: n5470_o = n5469_o;
    endcase
  assign n5471_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5472_o = n5471_o;
      13'b0100000000000: n5472_o = n5471_o;
      13'b0010000000000: n5472_o = n5471_o;
      13'b0001000000000: n5472_o = n5471_o;
      13'b0000100000000: n5472_o = n5471_o;
      13'b0000010000000: n5472_o = n5471_o;
      13'b0000001000000: n5472_o = n5471_o;
      13'b0000000100000: n5472_o = n5471_o;
      13'b0000000010000: n5472_o = n5471_o;
      13'b0000000001000: n5472_o = n5471_o;
      13'b0000000000100: n5472_o = n5471_o;
      13'b0000000000010: n5472_o = n5079_o;
      13'b0000000000001: n5472_o = n5471_o;
      default: n5472_o = n5471_o;
    endcase
  assign n5473_o = n2121_o[0];
  assign n5474_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5475_o = n1996_o ? n5473_o : n5474_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5476_o = n5475_o;
      13'b0100000000000: n5476_o = n5475_o;
      13'b0010000000000: n5476_o = n5352_o;
      13'b0001000000000: n5476_o = n5334_o;
      13'b0000100000000: n5476_o = n5312_o;
      13'b0000010000000: n5476_o = n5475_o;
      13'b0000001000000: n5476_o = n5475_o;
      13'b0000000100000: n5476_o = n5475_o;
      13'b0000000010000: n5476_o = n5475_o;
      13'b0000000001000: n5476_o = n5475_o;
      13'b0000000000100: n5476_o = n5475_o;
      13'b0000000000010: n5476_o = n5475_o;
      13'b0000000000001: n5476_o = n5475_o;
      default: n5476_o = n5475_o;
    endcase
  assign n5477_o = n2121_o[1];
  assign n5478_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5479_o = n1996_o ? n5477_o : n5478_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5480_o = n5479_o;
      13'b0100000000000: n5480_o = n5479_o;
      13'b0010000000000: n5480_o = n5479_o;
      13'b0001000000000: n5480_o = n5479_o;
      13'b0000100000000: n5480_o = n5479_o;
      13'b0000010000000: n5480_o = n5479_o;
      13'b0000001000000: n5480_o = n5479_o;
      13'b0000000100000: n5480_o = n5479_o;
      13'b0000000010000: n5480_o = n5479_o;
      13'b0000000001000: n5480_o = n5479_o;
      13'b0000000000100: n5480_o = n5479_o;
      13'b0000000000010: n5480_o = n5083_o;
      13'b0000000000001: n5480_o = n5479_o;
      default: n5480_o = n5479_o;
    endcase
  assign n5481_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5482_o = n5481_o;
      13'b0100000000000: n5482_o = n5481_o;
      13'b0010000000000: n5482_o = n5481_o;
      13'b0001000000000: n5482_o = n5481_o;
      13'b0000100000000: n5482_o = n5481_o;
      13'b0000010000000: n5482_o = n5481_o;
      13'b0000001000000: n5482_o = n5481_o;
      13'b0000000100000: n5482_o = n5481_o;
      13'b0000000010000: n5482_o = n5481_o;
      13'b0000000001000: n5482_o = n5481_o;
      13'b0000000000100: n5482_o = 1'b1;
      13'b0000000000010: n5482_o = 1'b1;
      13'b0000000000001: n5482_o = n5481_o;
      default: n5482_o = n5481_o;
    endcase
  assign n5483_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5484_o = n5483_o;
      13'b0100000000000: n5484_o = n5483_o;
      13'b0010000000000: n5484_o = n5483_o;
      13'b0001000000000: n5484_o = n5483_o;
      13'b0000100000000: n5484_o = n5483_o;
      13'b0000010000000: n5484_o = n5483_o;
      13'b0000001000000: n5484_o = n5483_o;
      13'b0000000100000: n5484_o = n5483_o;
      13'b0000000010000: n5484_o = n5483_o;
      13'b0000000001000: n5484_o = n5483_o;
      13'b0000000000100: n5484_o = n5483_o;
      13'b0000000000010: n5484_o = n5085_o;
      13'b0000000000001: n5484_o = n5483_o;
      default: n5484_o = n5483_o;
    endcase
  assign n5485_o = n1870_o[58:57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5486_o = n5485_o;
      13'b0100000000000: n5486_o = n5485_o;
      13'b0010000000000: n5486_o = n5354_o;
      13'b0001000000000: n5486_o = n5336_o;
      13'b0000100000000: n5486_o = n5485_o;
      13'b0000010000000: n5486_o = n5485_o;
      13'b0000001000000: n5486_o = n5485_o;
      13'b0000000100000: n5486_o = n5485_o;
      13'b0000000010000: n5486_o = n5485_o;
      13'b0000000001000: n5486_o = n5485_o;
      13'b0000000000100: n5486_o = n5485_o;
      13'b0000000000010: n5486_o = n5485_o;
      13'b0000000000001: n5486_o = n5485_o;
      default: n5486_o = n5485_o;
    endcase
  assign n5487_o = n1870_o[60:59];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5488_o = n5487_o;
      13'b0100000000000: n5488_o = n5487_o;
      13'b0010000000000: n5488_o = n5487_o;
      13'b0001000000000: n5488_o = n5487_o;
      13'b0000100000000: n5488_o = n5298_o;
      13'b0000010000000: n5488_o = n5487_o;
      13'b0000001000000: n5488_o = n5487_o;
      13'b0000000100000: n5488_o = n5487_o;
      13'b0000000010000: n5488_o = n5487_o;
      13'b0000000001000: n5488_o = n5487_o;
      13'b0000000000100: n5488_o = n5487_o;
      13'b0000000000010: n5488_o = n5487_o;
      13'b0000000000001: n5488_o = n5487_o;
      default: n5488_o = n5487_o;
    endcase
  assign n5489_o = n5423_o[0];
  assign n5490_o = n1976_o[0];
  assign n5491_o = n1870_o[65];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:17  */
  assign n5492_o = n1969_o ? n5490_o : n5491_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5493_o = n5489_o;
      13'b0100000000000: n5493_o = n5492_o;
      13'b0010000000000: n5493_o = n5492_o;
      13'b0001000000000: n5493_o = n5492_o;
      13'b0000100000000: n5493_o = n5492_o;
      13'b0000010000000: n5493_o = n5492_o;
      13'b0000001000000: n5493_o = n5492_o;
      13'b0000000100000: n5493_o = n5492_o;
      13'b0000000010000: n5493_o = n5492_o;
      13'b0000000001000: n5493_o = n5173_o;
      13'b0000000000100: n5493_o = n5492_o;
      13'b0000000000010: n5493_o = n5492_o;
      13'b0000000000001: n5493_o = n5492_o;
      default: n5493_o = n5492_o;
    endcase
  assign n5494_o = n5423_o[1];
  assign n5495_o = n1976_o[1];
  assign n5496_o = n1870_o[66];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1570:17  */
  assign n5497_o = n1969_o ? n5495_o : n5496_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5498_o = n5494_o;
      13'b0100000000000: n5498_o = n5497_o;
      13'b0010000000000: n5498_o = n5497_o;
      13'b0001000000000: n5498_o = n5497_o;
      13'b0000100000000: n5498_o = n5497_o;
      13'b0000010000000: n5498_o = n5497_o;
      13'b0000001000000: n5498_o = n5497_o;
      13'b0000000100000: n5498_o = n5497_o;
      13'b0000000010000: n5498_o = n5210_o;
      13'b0000000001000: n5498_o = n5497_o;
      13'b0000000000100: n5498_o = n5497_o;
      13'b0000000000010: n5498_o = n5497_o;
      13'b0000000000001: n5498_o = n5497_o;
      default: n5498_o = n5497_o;
    endcase
  assign n5499_o = n1870_o[74];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5500_o = n5499_o;
      13'b0100000000000: n5500_o = n5499_o;
      13'b0010000000000: n5500_o = n5499_o;
      13'b0001000000000: n5500_o = n5499_o;
      13'b0000100000000: n5500_o = n5499_o;
      13'b0000010000000: n5500_o = n5499_o;
      13'b0000001000000: n5500_o = n5499_o;
      13'b0000000100000: n5500_o = n5253_o;
      13'b0000000010000: n5500_o = n5499_o;
      13'b0000000001000: n5500_o = n5499_o;
      13'b0000000000100: n5500_o = n5499_o;
      13'b0000000000010: n5500_o = n5499_o;
      13'b0000000000001: n5500_o = n5499_o;
      default: n5500_o = n5499_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5502_o = 1'b0;
      13'b0100000000000: n5502_o = 1'b0;
      13'b0010000000000: n5502_o = 1'b0;
      13'b0001000000000: n5502_o = 1'b0;
      13'b0000100000000: n5502_o = 1'b0;
      13'b0000010000000: n5502_o = 1'b0;
      13'b0000001000000: n5502_o = 1'b0;
      13'b0000000100000: n5502_o = 1'b0;
      13'b0000000010000: n5502_o = 1'b0;
      13'b0000000001000: n5502_o = 1'b0;
      13'b0000000000100: n5502_o = 1'b1;
      13'b0000000000010: n5502_o = 1'b0;
      13'b0000000000001: n5502_o = 1'b0;
      default: n5502_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5504_o = 1'b0;
      13'b0100000000000: n5504_o = 1'b0;
      13'b0010000000000: n5504_o = 1'b0;
      13'b0001000000000: n5504_o = 1'b0;
      13'b0000100000000: n5504_o = 1'b0;
      13'b0000010000000: n5504_o = 1'b0;
      13'b0000001000000: n5504_o = 1'b0;
      13'b0000000100000: n5504_o = 1'b0;
      13'b0000000010000: n5504_o = 1'b0;
      13'b0000000001000: n5504_o = 1'b0;
      13'b0000000000100: n5504_o = 1'b0;
      13'b0000000000010: n5504_o = 1'b1;
      13'b0000000000001: n5504_o = 1'b0;
      default: n5504_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5506_o = n5425_o;
      13'b0100000000000: n5506_o = 2'b00;
      13'b0010000000000: n5506_o = 2'b00;
      13'b0001000000000: n5506_o = 2'b00;
      13'b0000100000000: n5506_o = 2'b00;
      13'b0000010000000: n5506_o = 2'b00;
      13'b0000001000000: n5506_o = 2'b00;
      13'b0000000100000: n5506_o = 2'b00;
      13'b0000000010000: n5506_o = 2'b00;
      13'b0000000001000: n5506_o = 2'b00;
      13'b0000000000100: n5506_o = 2'b00;
      13'b0000000000010: n5506_o = 2'b00;
      13'b0000000000001: n5506_o = 2'b00;
      default: n5506_o = 2'b00;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5508_o = 1'b0;
      13'b0100000000000: n5508_o = 1'b0;
      13'b0010000000000: n5508_o = 1'b0;
      13'b0001000000000: n5508_o = 1'b0;
      13'b0000100000000: n5508_o = 1'b0;
      13'b0000010000000: n5508_o = 1'b0;
      13'b0000001000000: n5508_o = 1'b0;
      13'b0000000100000: n5508_o = 1'b0;
      13'b0000000010000: n5508_o = n5212_o;
      13'b0000000001000: n5508_o = 1'b0;
      13'b0000000000100: n5508_o = 1'b1;
      13'b0000000000010: n5508_o = 1'b1;
      13'b0000000000001: n5508_o = 1'b0;
      default: n5508_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2455:65  */
  always @*
    case (n5432_o)
      13'b1000000000000: n5509_o = n5426_o;
      13'b0100000000000: n5509_o = n2139_o;
      13'b0010000000000: n5509_o = n5356_o;
      13'b0001000000000: n5509_o = n5338_o;
      13'b0000100000000: n5509_o = n5300_o;
      13'b0000010000000: n5509_o = n2139_o;
      13'b0000001000000: n5509_o = n2139_o;
      13'b0000000100000: n5509_o = n2139_o;
      13'b0000000010000: n5509_o = n2139_o;
      13'b0000000001000: n5509_o = n2139_o;
      13'b0000000000100: n5509_o = n5131_o;
      13'b0000000000010: n5509_o = n5087_o;
      13'b0000000000001: n5509_o = n2139_o;
      default: n5509_o = n2139_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5510_o = n4931_o ? n4990_o : n5433_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5511_o = n4931_o ? n4992_o : n5438_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5512_o = n4931_o ? n4993_o : n5439_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5513_o = n4931_o ? n2107_o : n5440_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5514_o = n4931_o ? n2110_o : n5441_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5515_o = n4931_o ? n4958_o : n5442_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5517_o = n4931_o ? n4996_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5519_o = n4931_o ? n4999_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5521_o = n4931_o ? 1'b0 : n5444_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5523_o = n4931_o ? 1'b0 : n5446_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5524_o = n4931_o ? n1867_o : n5447_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5525_o = n4931_o ? n2113_o : n5448_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5526_o = n4931_o ? n5002_o : n5451_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5528_o = n4931_o ? 1'b0 : n5453_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5530_o = n4931_o ? 1'b0 : n5456_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5532_o = n4931_o ? 1'b0 : n5458_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5533_o = n4931_o ? n5005_o : n5462_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5535_o = n4931_o ? 1'b0 : n5464_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5537_o = n4931_o ? n5008_o : 1'b0;
  assign n5538_o = {n5480_o, n5476_o};
  assign n5539_o = {n5488_o, n5486_o};
  assign n5540_o = {n5498_o, n5493_o};
  assign n5541_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5542_o = n4931_o ? n5541_o : n5466_o;
  assign n5543_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5544_o = n4931_o ? n5543_o : n5468_o;
  assign n5545_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5546_o = n4931_o ? n5545_o : n5470_o;
  assign n5547_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5548_o = n4931_o ? n5547_o : n5472_o;
  assign n5549_o = n5538_o[0];
  assign n5550_o = n2121_o[0];
  assign n5551_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5552_o = n1996_o ? n5550_o : n5551_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5553_o = n4931_o ? n5552_o : n5549_o;
  assign n5554_o = n5538_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5555_o = n4931_o ? n5013_o : n5554_o;
  assign n5556_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5557_o = n4931_o ? n5556_o : n5482_o;
  assign n5558_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5559_o = n4931_o ? n5558_o : n5484_o;
  assign n5560_o = n1870_o[60:57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5561_o = n4931_o ? n5560_o : n5539_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5562_o = n4931_o & n4944_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5563_o = n4931_o ? n1978_o : n5540_o;
  assign n5564_o = n1870_o[74];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5565_o = n4931_o ? n5564_o : n5500_o;
  assign n5566_o = {n5508_o, n5506_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5568_o = n4931_o ? 1'b0 : n5502_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5570_o = n4931_o ? 1'b0 : n5504_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5572_o = n4931_o ? 3'b000 : n5566_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2420:57  */
  assign n5573_o = n4931_o ? n5015_o : n5509_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2402:49  */
  assign n5575_o = n3568_o == 3'b111;
  assign n5576_o = {n5575_o, n4930_o, n4820_o, n4033_o, n3893_o, n3786_o, n3687_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5577_o = n5510_o;
      7'b0100000: n5577_o = make_berr;
      7'b0010000: n5577_o = make_berr;
      7'b0001000: n5577_o = make_berr;
      7'b0000100: n5577_o = make_berr;
      7'b0000010: n5577_o = n3767_o;
      7'b0000001: n5577_o = n3598_o;
      default: n5577_o = make_berr;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5578_o = n5511_o;
      7'b0100000: n5578_o = n4910_o;
      7'b0010000: n5578_o = n4740_o;
      7'b0001000: n5578_o = n3938_o;
      7'b0000100: n5578_o = n3815_o;
      7'b0000010: n5578_o = n3715_o;
      7'b0000001: n5578_o = n3607_o;
      default: n5578_o = n1882_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5579_o = n5512_o;
      7'b0100000: n5579_o = n1985_o;
      7'b0010000: n5579_o = n4741_o;
      7'b0001000: n5579_o = n3936_o;
      7'b0000100: n5579_o = n1985_o;
      7'b0000010: n5579_o = n1985_o;
      7'b0000001: n5579_o = n1985_o;
      default: n5579_o = n1985_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5580_o = n5513_o;
      7'b0100000: n5580_o = n2107_o;
      7'b0010000: n5580_o = n2107_o;
      7'b0001000: n5580_o = n2107_o;
      7'b0000100: n5580_o = n2107_o;
      7'b0000010: n5580_o = n2107_o;
      7'b0000001: n5580_o = n2107_o;
      default: n5580_o = n2107_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5581_o = n5514_o;
      7'b0100000: n5581_o = n2110_o;
      7'b0010000: n5581_o = n2110_o;
      7'b0001000: n5581_o = n2110_o;
      7'b0000100: n5581_o = n2110_o;
      7'b0000010: n5581_o = n2110_o;
      7'b0000001: n5581_o = n2110_o;
      default: n5581_o = n2110_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5583_o = 1'b0;
      7'b0100000: n5583_o = n4912_o;
      7'b0010000: n5583_o = n4743_o;
      7'b0001000: n5583_o = n4014_o;
      7'b0000100: n5583_o = n3877_o;
      7'b0000010: n5583_o = n3770_o;
      7'b0000001: n5583_o = n3663_o;
      default: n5583_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5584_o = n5515_o;
      7'b0100000: n5584_o = n1974_o;
      7'b0010000: n5584_o = n4744_o;
      7'b0001000: n5584_o = n1974_o;
      7'b0000100: n5584_o = n1974_o;
      7'b0000010: n5584_o = n1974_o;
      7'b0000001: n5584_o = n1974_o;
      default: n5584_o = n1974_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5586_o = n5517_o;
      7'b0100000: n5586_o = 1'b0;
      7'b0010000: n5586_o = 1'b0;
      7'b0001000: n5586_o = 1'b0;
      7'b0000100: n5586_o = 1'b0;
      7'b0000010: n5586_o = 1'b0;
      7'b0000001: n5586_o = 1'b0;
      default: n5586_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5588_o = 1'b0;
      7'b0100000: n5588_o = n4914_o;
      7'b0010000: n5588_o = 1'b0;
      7'b0001000: n5588_o = 1'b0;
      7'b0000100: n5588_o = 1'b0;
      7'b0000010: n5588_o = 1'b0;
      7'b0000001: n5588_o = 1'b0;
      default: n5588_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5590_o = n5519_o;
      7'b0100000: n5590_o = 1'b0;
      7'b0010000: n5590_o = n4745_o;
      7'b0001000: n5590_o = 1'b0;
      7'b0000100: n5590_o = 1'b0;
      7'b0000010: n5590_o = 1'b0;
      7'b0000001: n5590_o = 1'b0;
      default: n5590_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5592_o = n5521_o;
      7'b0100000: n5592_o = n4916_o;
      7'b0010000: n5592_o = n4747_o;
      7'b0001000: n5592_o = 1'b0;
      7'b0000100: n5592_o = 1'b0;
      7'b0000010: n5592_o = 1'b0;
      7'b0000001: n5592_o = 1'b0;
      default: n5592_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5594_o = n5523_o;
      7'b0100000: n5594_o = n4918_o;
      7'b0010000: n5594_o = n4748_o;
      7'b0001000: n5594_o = n4016_o;
      7'b0000100: n5594_o = n3878_o;
      7'b0000010: n5594_o = 1'b0;
      7'b0000001: n5594_o = n3665_o;
      default: n5594_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5596_o = 1'b0;
      7'b0100000: n5596_o = 1'b0;
      7'b0010000: n5596_o = n4750_o;
      7'b0001000: n5596_o = 1'b0;
      7'b0000100: n5596_o = 1'b0;
      7'b0000010: n5596_o = 1'b0;
      7'b0000001: n5596_o = 1'b0;
      default: n5596_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5598_o = 1'b0;
      7'b0100000: n5598_o = 1'b0;
      7'b0010000: n5598_o = n4752_o;
      7'b0001000: n5598_o = 1'b0;
      7'b0000100: n5598_o = 1'b0;
      7'b0000010: n5598_o = 1'b0;
      7'b0000001: n5598_o = 1'b0;
      default: n5598_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5600_o = 1'b0;
      7'b0100000: n5600_o = 1'b0;
      7'b0010000: n5600_o = n4754_o;
      7'b0001000: n5600_o = 1'b0;
      7'b0000100: n5600_o = 1'b0;
      7'b0000010: n5600_o = 1'b0;
      7'b0000001: n5600_o = 1'b0;
      default: n5600_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5601_o = n5524_o;
      7'b0100000: n5601_o = n1867_o;
      7'b0010000: n5601_o = n1867_o;
      7'b0001000: n5601_o = n1867_o;
      7'b0000100: n5601_o = n1867_o;
      7'b0000010: n5601_o = n1867_o;
      7'b0000001: n5601_o = n1867_o;
      default: n5601_o = n1867_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5603_o = 1'b0;
      7'b0100000: n5603_o = 1'b0;
      7'b0010000: n5603_o = n4756_o;
      7'b0001000: n5603_o = 1'b0;
      7'b0000100: n5603_o = 1'b0;
      7'b0000010: n5603_o = 1'b0;
      7'b0000001: n5603_o = 1'b0;
      default: n5603_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5604_o = n5525_o;
      7'b0100000: n5604_o = n2113_o;
      7'b0010000: n5604_o = n2113_o;
      7'b0001000: n5604_o = n2113_o;
      7'b0000100: n5604_o = n2113_o;
      7'b0000010: n5604_o = n2113_o;
      7'b0000001: n5604_o = n2113_o;
      default: n5604_o = n2113_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5606_o = n5526_o;
      7'b0100000: n5606_o = n4920_o;
      7'b0010000: n5606_o = n4757_o;
      7'b0001000: n5606_o = n4017_o;
      7'b0000100: n5606_o = n3879_o;
      7'b0000010: n5606_o = n3772_o;
      7'b0000001: n5606_o = n3668_o;
      default: n5606_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5608_o = n5528_o;
      7'b0100000: n5608_o = 1'b0;
      7'b0010000: n5608_o = 1'b0;
      7'b0001000: n5608_o = n4019_o;
      7'b0000100: n5608_o = 1'b0;
      7'b0000010: n5608_o = 1'b0;
      7'b0000001: n5608_o = n3670_o;
      default: n5608_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5610_o = n5530_o;
      7'b0100000: n5610_o = 1'b0;
      7'b0010000: n5610_o = 1'b0;
      7'b0001000: n5610_o = 1'b0;
      7'b0000100: n5610_o = 1'b0;
      7'b0000010: n5610_o = 1'b0;
      7'b0000001: n5610_o = 1'b0;
      default: n5610_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5612_o = n5532_o;
      7'b0100000: n5612_o = 1'b0;
      7'b0010000: n5612_o = 1'b0;
      7'b0001000: n5612_o = 1'b0;
      7'b0000100: n5612_o = 1'b0;
      7'b0000010: n5612_o = 1'b0;
      7'b0000001: n5612_o = 1'b0;
      default: n5612_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5614_o = n5533_o;
      7'b0100000: n5614_o = n4922_o;
      7'b0010000: n5614_o = n4758_o;
      7'b0001000: n5614_o = n4020_o;
      7'b0000100: n5614_o = n3880_o;
      7'b0000010: n5614_o = n3774_o;
      7'b0000001: n5614_o = n3672_o;
      default: n5614_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5616_o = n5535_o;
      7'b0100000: n5616_o = 1'b0;
      7'b0010000: n5616_o = 1'b0;
      7'b0001000: n5616_o = 1'b0;
      7'b0000100: n5616_o = 1'b0;
      7'b0000010: n5616_o = 1'b0;
      7'b0000001: n5616_o = 1'b0;
      default: n5616_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5618_o = n5537_o;
      7'b0100000: n5618_o = n4924_o;
      7'b0010000: n5618_o = n4760_o;
      7'b0001000: n5618_o = n4021_o;
      7'b0000100: n5618_o = n3881_o;
      7'b0000010: n5618_o = n3776_o;
      7'b0000001: n5618_o = n3674_o;
      default: n5618_o = 1'b0;
    endcase
  assign n5619_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5620_o = n5542_o;
      7'b0100000: n5620_o = n5619_o;
      7'b0010000: n5620_o = n4762_o;
      7'b0001000: n5620_o = n5619_o;
      7'b0000100: n5620_o = n5619_o;
      7'b0000010: n5620_o = n5619_o;
      7'b0000001: n5620_o = n5619_o;
      default: n5620_o = n5619_o;
    endcase
  assign n5621_o = n1870_o[20];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5622_o = n5621_o;
      7'b0100000: n5622_o = n5621_o;
      7'b0010000: n5622_o = n4764_o;
      7'b0001000: n5622_o = n5621_o;
      7'b0000100: n5622_o = n5621_o;
      7'b0000010: n5622_o = n5621_o;
      7'b0000001: n5622_o = n5621_o;
      default: n5622_o = n5621_o;
    endcase
  assign n5623_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5624_o = n5544_o;
      7'b0100000: n5624_o = n5623_o;
      7'b0010000: n5624_o = n4766_o;
      7'b0001000: n5624_o = n5623_o;
      7'b0000100: n5624_o = n5623_o;
      7'b0000010: n5624_o = n5623_o;
      7'b0000001: n5624_o = n5623_o;
      default: n5624_o = n5623_o;
    endcase
  assign n5625_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5626_o = n5546_o;
      7'b0100000: n5626_o = n5625_o;
      7'b0010000: n5626_o = n4767_o;
      7'b0001000: n5626_o = n5625_o;
      7'b0000100: n5626_o = n5625_o;
      7'b0000010: n5626_o = n5625_o;
      7'b0000001: n5626_o = n5625_o;
      default: n5626_o = n5625_o;
    endcase
  assign n5627_o = n1870_o[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5628_o = n5627_o;
      7'b0100000: n5628_o = n5627_o;
      7'b0010000: n5628_o = n4769_o;
      7'b0001000: n5628_o = n5627_o;
      7'b0000100: n5628_o = n5627_o;
      7'b0000010: n5628_o = n5627_o;
      7'b0000001: n5628_o = n5627_o;
      default: n5628_o = n5627_o;
    endcase
  assign n5629_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5630_o = n5629_o;
      7'b0100000: n5630_o = n5629_o;
      7'b0010000: n5630_o = n4771_o;
      7'b0001000: n5630_o = n5629_o;
      7'b0000100: n5630_o = n5629_o;
      7'b0000010: n5630_o = n5629_o;
      7'b0000001: n5630_o = n5629_o;
      default: n5630_o = n5629_o;
    endcase
  assign n5631_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5632_o = n5631_o;
      7'b0100000: n5632_o = n5631_o;
      7'b0010000: n5632_o = n4772_o;
      7'b0001000: n5632_o = n5631_o;
      7'b0000100: n5632_o = n5631_o;
      7'b0000010: n5632_o = n5631_o;
      7'b0000001: n5632_o = n5631_o;
      default: n5632_o = n5631_o;
    endcase
  assign n5633_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5634_o = n5548_o;
      7'b0100000: n5634_o = n5633_o;
      7'b0010000: n5634_o = n4774_o;
      7'b0001000: n5634_o = n5633_o;
      7'b0000100: n5634_o = n5633_o;
      7'b0000010: n5634_o = n5633_o;
      7'b0000001: n5634_o = n5633_o;
      default: n5634_o = n5633_o;
    endcase
  assign n5635_o = n2121_o[0];
  assign n5636_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5637_o = n1996_o ? n5635_o : n5636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5638_o = n5553_o;
      7'b0100000: n5638_o = n5637_o;
      7'b0010000: n5638_o = n5637_o;
      7'b0001000: n5638_o = n5637_o;
      7'b0000100: n5638_o = n5637_o;
      7'b0000010: n5638_o = n5637_o;
      7'b0000001: n5638_o = n5637_o;
      default: n5638_o = n5637_o;
    endcase
  assign n5639_o = n2121_o[1];
  assign n5640_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n5641_o = n1996_o ? n5639_o : n5640_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5642_o = n5555_o;
      7'b0100000: n5642_o = n5641_o;
      7'b0010000: n5642_o = n4778_o;
      7'b0001000: n5642_o = n5641_o;
      7'b0000100: n5642_o = n5641_o;
      7'b0000010: n5642_o = n5641_o;
      7'b0000001: n5642_o = n5641_o;
      default: n5642_o = n5641_o;
    endcase
  assign n5643_o = n1870_o[48];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5644_o = n5643_o;
      7'b0100000: n5644_o = n5643_o;
      7'b0010000: n5644_o = n4781_o;
      7'b0001000: n5644_o = n5643_o;
      7'b0000100: n5644_o = n5643_o;
      7'b0000010: n5644_o = n5643_o;
      7'b0000001: n5644_o = n5643_o;
      default: n5644_o = n5643_o;
    endcase
  assign n5645_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5646_o = n5557_o;
      7'b0100000: n5646_o = n5645_o;
      7'b0010000: n5646_o = n4783_o;
      7'b0001000: n5646_o = n5645_o;
      7'b0000100: n5646_o = n5645_o;
      7'b0000010: n5646_o = n5645_o;
      7'b0000001: n5646_o = n5645_o;
      default: n5646_o = n5645_o;
    endcase
  assign n5647_o = n3922_o[0];
  assign n5648_o = n1870_o[51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5649_o = n5648_o;
      7'b0100000: n5649_o = n5648_o;
      7'b0010000: n5649_o = n5648_o;
      7'b0001000: n5649_o = n5647_o;
      7'b0000100: n5649_o = n3813_o;
      7'b0000010: n5649_o = n5648_o;
      7'b0000001: n5649_o = n5648_o;
      default: n5649_o = n5648_o;
    endcase
  assign n5650_o = n3922_o[1];
  assign n5651_o = n1870_o[52];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5652_o = n5651_o;
      7'b0100000: n5652_o = n5651_o;
      7'b0010000: n5652_o = n5651_o;
      7'b0001000: n5652_o = n5650_o;
      7'b0000100: n5652_o = n5651_o;
      7'b0000010: n5652_o = n5651_o;
      7'b0000001: n5652_o = n5651_o;
      default: n5652_o = n5651_o;
    endcase
  assign n5653_o = n1870_o[53];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5654_o = n5653_o;
      7'b0100000: n5654_o = n5653_o;
      7'b0010000: n5654_o = n5653_o;
      7'b0001000: n5654_o = n4025_o;
      7'b0000100: n5654_o = n5653_o;
      7'b0000010: n5654_o = n5653_o;
      7'b0000001: n5654_o = n5653_o;
      default: n5654_o = n5653_o;
    endcase
  assign n5655_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5656_o = n5655_o;
      7'b0100000: n5656_o = n5655_o;
      7'b0010000: n5656_o = n4786_o;
      7'b0001000: n5656_o = n5655_o;
      7'b0000100: n5656_o = n3885_o;
      7'b0000010: n5656_o = n3778_o;
      7'b0000001: n5656_o = n3676_o;
      default: n5656_o = n5655_o;
    endcase
  assign n5657_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5658_o = n5559_o;
      7'b0100000: n5658_o = n5657_o;
      7'b0010000: n5658_o = n4788_o;
      7'b0001000: n5658_o = n5657_o;
      7'b0000100: n5658_o = n5657_o;
      7'b0000010: n5658_o = n5657_o;
      7'b0000001: n5658_o = n5657_o;
      default: n5658_o = n5657_o;
    endcase
  assign n5659_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5660_o = n5659_o;
      7'b0100000: n5660_o = n5659_o;
      7'b0010000: n5660_o = n4791_o;
      7'b0001000: n5660_o = n5659_o;
      7'b0000100: n5660_o = n3887_o;
      7'b0000010: n5660_o = n5659_o;
      7'b0000001: n5660_o = n3678_o;
      default: n5660_o = n5659_o;
    endcase
  assign n5661_o = n1870_o[60:57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5662_o = n5561_o;
      7'b0100000: n5662_o = n5661_o;
      7'b0010000: n5662_o = n5661_o;
      7'b0001000: n5662_o = n5661_o;
      7'b0000100: n5662_o = n5661_o;
      7'b0000010: n5662_o = n5661_o;
      7'b0000001: n5662_o = n5661_o;
      default: n5662_o = n5661_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5663_o = n5014_o;
      7'b0100000: n5663_o = n2137_o;
      7'b0010000: n5663_o = n2137_o;
      7'b0001000: n5663_o = n2137_o;
      7'b0000100: n5663_o = n2137_o;
      7'b0000010: n5663_o = n2137_o;
      7'b0000001: n5663_o = n2137_o;
      default: n5663_o = n2137_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5664_o = n5563_o;
      7'b0100000: n5664_o = n1978_o;
      7'b0010000: n5664_o = n1978_o;
      7'b0001000: n5664_o = n1978_o;
      7'b0000100: n5664_o = n1978_o;
      7'b0000010: n5664_o = n1978_o;
      7'b0000001: n5664_o = n1978_o;
      default: n5664_o = n1978_o;
    endcase
  assign n5665_o = n1870_o[67];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5666_o = n5665_o;
      7'b0100000: n5666_o = n5665_o;
      7'b0010000: n5666_o = n4793_o;
      7'b0001000: n5666_o = n5665_o;
      7'b0000100: n5666_o = n5665_o;
      7'b0000010: n5666_o = n5665_o;
      7'b0000001: n5666_o = n5665_o;
      default: n5666_o = n5665_o;
    endcase
  assign n5667_o = n1870_o[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5668_o = n5667_o;
      7'b0100000: n5668_o = n5667_o;
      7'b0010000: n5668_o = n4795_o;
      7'b0001000: n5668_o = n5667_o;
      7'b0000100: n5668_o = n5667_o;
      7'b0000010: n5668_o = n5667_o;
      7'b0000001: n5668_o = n5667_o;
      default: n5668_o = n5667_o;
    endcase
  assign n5669_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5670_o = n5669_o;
      7'b0100000: n5670_o = n5669_o;
      7'b0010000: n5670_o = n4796_o;
      7'b0001000: n5670_o = n5669_o;
      7'b0000100: n5670_o = n5669_o;
      7'b0000010: n5670_o = n5669_o;
      7'b0000001: n5670_o = n5669_o;
      default: n5670_o = n5669_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5671_o = n2130_o;
      7'b0100000: n5671_o = n2130_o;
      7'b0010000: n5671_o = n4797_o;
      7'b0001000: n5671_o = n2130_o;
      7'b0000100: n5671_o = n2130_o;
      7'b0000010: n5671_o = n2130_o;
      7'b0000001: n5671_o = n2130_o;
      default: n5671_o = n2130_o;
    endcase
  assign n5672_o = n1870_o[74];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5673_o = n5565_o;
      7'b0100000: n5673_o = n5672_o;
      7'b0010000: n5673_o = n5672_o;
      7'b0001000: n5673_o = n5672_o;
      7'b0000100: n5673_o = n5672_o;
      7'b0000010: n5673_o = n5672_o;
      7'b0000001: n5673_o = n5672_o;
      default: n5673_o = n5672_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5675_o = n5568_o;
      7'b0100000: n5675_o = n4926_o;
      7'b0010000: n5675_o = n4799_o;
      7'b0001000: n5675_o = 1'b0;
      7'b0000100: n5675_o = 1'b0;
      7'b0000010: n5675_o = 1'b0;
      7'b0000001: n5675_o = 1'b0;
      default: n5675_o = 1'b0;
    endcase
  assign n5676_o = n3681_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5678_o = 1'b0;
      7'b0100000: n5678_o = 1'b0;
      7'b0010000: n5678_o = 1'b0;
      7'b0001000: n5678_o = 1'b0;
      7'b0000100: n5678_o = 1'b0;
      7'b0000010: n5678_o = n3780_o;
      7'b0000001: n5678_o = n5676_o;
      default: n5678_o = 1'b0;
    endcase
  assign n5679_o = n3681_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5681_o = n5570_o;
      7'b0100000: n5681_o = 1'b0;
      7'b0010000: n5681_o = n4801_o;
      7'b0001000: n5681_o = 1'b0;
      7'b0000100: n5681_o = n3889_o;
      7'b0000010: n5681_o = 1'b0;
      7'b0000001: n5681_o = n5679_o;
      default: n5681_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5683_o = 1'b0;
      7'b0100000: n5683_o = 1'b0;
      7'b0010000: n5683_o = 1'b0;
      7'b0001000: n5683_o = 1'b0;
      7'b0000100: n5683_o = 1'b0;
      7'b0000010: n5683_o = n3782_o;
      7'b0000001: n5683_o = 1'b0;
      default: n5683_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5685_o = 1'b0;
      7'b0100000: n5685_o = 1'b0;
      7'b0010000: n5685_o = 1'b0;
      7'b0001000: n5685_o = n4027_o;
      7'b0000100: n5685_o = 1'b0;
      7'b0000010: n5685_o = 1'b0;
      7'b0000001: n5685_o = 1'b0;
      default: n5685_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5687_o = 1'b0;
      7'b0100000: n5687_o = 1'b0;
      7'b0010000: n5687_o = n4803_o;
      7'b0001000: n5687_o = 1'b0;
      7'b0000100: n5687_o = 1'b0;
      7'b0000010: n5687_o = 1'b0;
      7'b0000001: n5687_o = 1'b0;
      default: n5687_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5689_o = 1'b0;
      7'b0100000: n5689_o = 1'b0;
      7'b0010000: n5689_o = n4805_o;
      7'b0001000: n5689_o = 1'b0;
      7'b0000100: n5689_o = 1'b0;
      7'b0000010: n5689_o = 1'b0;
      7'b0000001: n5689_o = 1'b0;
      default: n5689_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5691_o = 1'b0;
      7'b0100000: n5691_o = 1'b0;
      7'b0010000: n5691_o = n4807_o;
      7'b0001000: n5691_o = 1'b0;
      7'b0000100: n5691_o = 1'b0;
      7'b0000010: n5691_o = 1'b0;
      7'b0000001: n5691_o = 1'b0;
      default: n5691_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5693_o = 1'b0;
      7'b0100000: n5693_o = 1'b0;
      7'b0010000: n5693_o = 1'b0;
      7'b0001000: n5693_o = n4029_o;
      7'b0000100: n5693_o = 1'b0;
      7'b0000010: n5693_o = 1'b0;
      7'b0000001: n5693_o = 1'b0;
      default: n5693_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5695_o = 1'b0;
      7'b0100000: n5695_o = 1'b0;
      7'b0010000: n5695_o = n4809_o;
      7'b0001000: n5695_o = 1'b0;
      7'b0000100: n5695_o = 1'b0;
      7'b0000010: n5695_o = 1'b0;
      7'b0000001: n5695_o = n3683_o;
      default: n5695_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5697_o = 1'b0;
      7'b0100000: n5697_o = 1'b0;
      7'b0010000: n5697_o = n4811_o;
      7'b0001000: n5697_o = 1'b0;
      7'b0000100: n5697_o = 1'b0;
      7'b0000010: n5697_o = 1'b0;
      7'b0000001: n5697_o = 1'b0;
      default: n5697_o = 1'b0;
    endcase
  assign n5698_o = n5572_o[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5700_o = n5698_o;
      7'b0100000: n5700_o = 2'b00;
      7'b0010000: n5700_o = 2'b00;
      7'b0001000: n5700_o = 2'b00;
      7'b0000100: n5700_o = 2'b00;
      7'b0000010: n5700_o = 2'b00;
      7'b0000001: n5700_o = 2'b00;
      default: n5700_o = 2'b00;
    endcase
  assign n5701_o = n5572_o[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5703_o = n5701_o;
      7'b0100000: n5703_o = n4928_o;
      7'b0010000: n5703_o = n4812_o;
      7'b0001000: n5703_o = n4031_o;
      7'b0000100: n5703_o = n3891_o;
      7'b0000010: n5703_o = n3784_o;
      7'b0000001: n5703_o = n3685_o;
      default: n5703_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5705_o = 1'b0;
      7'b0100000: n5705_o = 1'b0;
      7'b0010000: n5705_o = n4814_o;
      7'b0001000: n5705_o = 1'b0;
      7'b0000100: n5705_o = 1'b0;
      7'b0000010: n5705_o = 1'b0;
      7'b0000001: n5705_o = 1'b0;
      default: n5705_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2031:41  */
  always @*
    case (n5576_o)
      7'b1000000: n5706_o = n5573_o;
      7'b0100000: n5706_o = n2139_o;
      7'b0010000: n5706_o = n4815_o;
      7'b0001000: n5706_o = n2139_o;
      7'b0000100: n5706_o = n2139_o;
      7'b0000010: n5706_o = n2139_o;
      7'b0000001: n5706_o = n2139_o;
      default: n5706_o = n2139_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5707_o = n3311_o ? make_berr : n5577_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5708_o = n3311_o ? n3538_o : n5578_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5709_o = n3311_o ? n3539_o : n5579_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5710_o = n3311_o ? n2107_o : n5580_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5711_o = n3311_o ? n2110_o : n5581_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5713_o = n3311_o ? 1'b0 : n5583_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5714_o = n3311_o ? n1974_o : n5584_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5716_o = n3311_o ? 1'b0 : n5586_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5718_o = n3311_o ? 1'b0 : n5588_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5719_o = n3311_o ? n3541_o : n5590_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5720_o = n3311_o ? n3543_o : n5592_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5721_o = n3311_o ? n3544_o : n5594_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5723_o = n3311_o ? 1'b0 : n5596_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5725_o = n3311_o ? n3546_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5727_o = n3311_o ? 1'b0 : n5598_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5728_o = n3311_o ? n3547_o : n5600_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5729_o = n3311_o ? n1867_o : n5601_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5731_o = n3311_o ? 1'b0 : n5603_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5732_o = n3311_o ? n3548_o : n5604_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5733_o = n3311_o ? n3549_o : n5606_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5735_o = n3311_o ? 1'b0 : n5608_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5737_o = n3311_o ? 1'b0 : n5610_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5739_o = n3311_o ? 1'b0 : n5612_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5740_o = n3311_o ? n3550_o : n5614_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5742_o = n3311_o ? 1'b0 : n5616_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5743_o = n3311_o ? n3551_o : n5618_o;
  assign n5744_o = {n5646_o, n5644_o, n5642_o, n5638_o};
  assign n5745_o = {n5662_o, n5660_o, n5658_o, n5656_o, n5654_o, n5652_o, n5649_o};
  assign n5746_o = {n5666_o, n5664_o, n5663_o};
  assign n5747_o = {n5673_o, n5671_o};
  assign n5748_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5749_o = n3311_o ? n5748_o : n5620_o;
  assign n5750_o = n1870_o[20];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5751_o = n3311_o ? n5750_o : n5622_o;
  assign n5752_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5753_o = n3311_o ? n5752_o : n5624_o;
  assign n5754_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5755_o = n3311_o ? n5754_o : n5626_o;
  assign n5756_o = n1870_o[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5757_o = n3311_o ? n5756_o : n5628_o;
  assign n5758_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5759_o = n3311_o ? n5758_o : n5630_o;
  assign n5760_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5761_o = n3311_o ? n5760_o : n5632_o;
  assign n5762_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5763_o = n3311_o ? n3553_o : n5762_o;
  assign n5764_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5765_o = n3311_o ? n5764_o : n5634_o;
  assign n5766_o = n5744_o[2:0];
  assign n5767_o = n1870_o[48];
  assign n5768_o = {n5767_o, n2125_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5769_o = n3311_o ? n5768_o : n5766_o;
  assign n5770_o = n5744_o[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5771_o = n3311_o ? n3555_o : n5770_o;
  assign n5772_o = n5745_o[4:0];
  assign n5773_o = n1870_o[55:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5774_o = n3311_o ? n5773_o : n5772_o;
  assign n5775_o = n5745_o[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5776_o = n3311_o ? n3557_o : n5775_o;
  assign n5777_o = n5745_o[9:6];
  assign n5778_o = n1870_o[60:57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5779_o = n3311_o ? n5778_o : n5777_o;
  assign n5780_o = n1870_o[67];
  assign n5781_o = {n5780_o, n1978_o, n2137_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5782_o = n3311_o ? n5781_o : n5746_o;
  assign n5783_o = n1870_o[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5784_o = n3311_o ? n5783_o : n5668_o;
  assign n5785_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5786_o = n3311_o ? n5785_o : n5670_o;
  assign n5787_o = n1870_o[74];
  assign n5788_o = {n5787_o, n2130_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5789_o = n3311_o ? n5788_o : n5747_o;
  assign n5790_o = {n5681_o, n5678_o};
  assign n5791_o = {n5685_o, n5683_o};
  assign n5792_o = {n5703_o, n5700_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5793_o = n3311_o ? n3559_o : n5675_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5795_o = n3311_o ? 2'b00 : n5790_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5797_o = n3311_o ? 2'b00 : n5791_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5798_o = n3311_o ? n3561_o : n5687_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5800_o = n3311_o ? 1'b0 : n5689_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5802_o = n3311_o ? 1'b0 : n5691_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5804_o = n3311_o ? 1'b0 : n5693_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5806_o = n3311_o ? 1'b0 : n5695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5808_o = n3311_o ? 1'b0 : n5697_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5810_o = n3311_o ? n3563_o : 1'b0;
  assign n5811_o = n5792_o[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5813_o = n3311_o ? 2'b00 : n5811_o;
  assign n5814_o = n5792_o[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5815_o = n3311_o ? n3565_o : n5814_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5816_o = n3311_o ? n3567_o : n5705_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1953:33  */
  assign n5817_o = n3311_o ? n2139_o : n5706_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1952:25  */
  assign n5819_o = n2140_o == 4'b0100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:50  */
  assign n5820_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:62  */
  assign n5822_o = n5820_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:58  */
  assign n5823_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:70  */
  assign n5825_o = n5823_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2633:57  */
  assign n5829_o = decodeopc ? 1'b1 : 1'b0;
  assign n5830_o = n1870_o[53];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n5831_o = n6026_o ? 1'b1 : n5830_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2633:57  */
  assign n5833_o = decodeopc ? 7'b0011001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:61  */
  assign n5834_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:73  */
  assign n5836_o = n5834_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:91  */
  assign n5837_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:103  */
  assign n5839_o = n5837_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:118  */
  assign n5840_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:130  */
  assign n5842_o = n5840_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:109  */
  assign n5843_o = n5839_o | n5842_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:80  */
  assign n5844_o = n5836_o & n5843_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2639:63  */
  assign n5845_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2640:74  */
  assign n5846_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2640:86  */
  assign n5848_o = n5846_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2642:90  */
  assign n5849_o = opcode[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5851_o = n5930_o ? 1'b1 : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2641:73  */
  assign n5852_o = decodeopc & n5849_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5854_o = n5935_o ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2648:73  */
  assign n5856_o = decodeopc ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2640:65  */
  assign n5857_o = n5848_o ? n1985_o : n5856_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2640:65  */
  assign n5858_o = n5848_o & n5852_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2640:65  */
  assign n5859_o = n5848_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2652:99  */
  assign n5860_o = ~decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2652:86  */
  assign n5861_o = exe_condition & n5860_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2652:65  */
  assign n5864_o = n5861_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2652:65  */
  assign n5867_o = n5861_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5868_o = n5921_o ? n5857_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2639:57  */
  assign n5871_o = n5845_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2639:57  */
  assign n5873_o = n5845_o ? n5864_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2639:57  */
  assign n5875_o = n5845_o ? n5867_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2639:57  */
  assign n5876_o = n5845_o & n5858_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2639:57  */
  assign n5877_o = n5845_o & n5859_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:62  */
  assign n5878_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:74  */
  assign n5880_o = n5878_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:91  */
  assign n5881_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:103  */
  assign n5883_o = n5881_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:82  */
  assign n5884_o = n5880_o | n5883_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2665:63  */
  assign n5886_o = cpu[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2665:80  */
  assign n5888_o = state == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2665:71  */
  assign n5889_o = n5886_o & n5888_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2665:99  */
  assign n5890_o = ~addrvalue;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2665:86  */
  assign n5891_o = n5889_o & n5890_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5893_o = n5900_o ? 1'b1 : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2668:66  */
  assign n5894_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2668:78  */
  assign n5896_o = n5894_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2668:57  */
  assign n5899_o = n5896_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5900_o = n5884_o & n5891_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5902_o = n5884_o ? 2'b00 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5905_o = n5884_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5908_o = n5884_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5911_o = n5884_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5914_o = n5884_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5916_o = n5884_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2660:49  */
  assign n5918_o = n5884_o ? n5899_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5919_o = n5844_o ? make_berr : n5893_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5920_o = n5844_o ? n1882_o : n5902_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5921_o = n5844_o & n5845_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5923_o = n5844_o ? 1'b0 : n5905_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5924_o = n5844_o ? n5871_o : n5908_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5926_o = n5844_o ? n5873_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5927_o = n5844_o ? n5875_o : n5911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5929_o = n5844_o ? 1'b0 : n5914_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5930_o = n5844_o & n5876_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5932_o = n5844_o ? 1'b0 : n5916_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5934_o = n5844_o ? 1'b0 : n5918_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2638:49  */
  assign n5935_o = n5844_o & n5877_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5936_o = n5825_o ? make_berr : n5919_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5937_o = n5825_o ? n1882_o : n5920_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5938_o = n5825_o ? n1985_o : n5868_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5940_o = n5825_o ? n5829_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5942_o = n5825_o ? 1'b0 : n5923_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5944_o = n5825_o ? 1'b0 : n5924_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5946_o = n5825_o ? 1'b0 : n5926_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5948_o = n5825_o ? 1'b0 : n5927_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5950_o = n5825_o ? 1'b0 : n5929_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5952_o = n5825_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5953_o = n5825_o ? n2130_o : n5851_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5955_o = n5825_o ? 1'b0 : n5932_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5957_o = n5825_o ? 1'b0 : n5934_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2632:49  */
  assign n5958_o = n5825_o ? n5833_o : n5854_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:58  */
  assign n5959_o = opcode[7:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:70  */
  assign n5961_o = n5959_o != 5'b00001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2677:59  */
  assign n5962_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2677:71  */
  assign n5964_o = n5962_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2677:88  */
  assign n5965_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2677:100  */
  assign n5967_o = n5965_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2677:79  */
  assign n5968_o = n5964_o | n5967_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:80  */
  assign n5969_o = n5961_o & n5968_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2679:66  */
  assign n5970_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2679:78  */
  assign n5972_o = n5970_o == 3'b001;
  assign n5974_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n5975_o = n6002_o ? 1'b1 : n5974_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2682:66  */
  assign n5976_o = opcode[8];
  assign n5978_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n5979_o = n6004_o ? 1'b1 : n5978_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2689:66  */
  assign n5983_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2689:78  */
  assign n5985_o = n5983_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2689:57  */
  assign n5988_o = n5985_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n5991_o = n5969_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n5994_o = n5969_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n5997_o = n5969_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n6000_o = n5969_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n6002_o = n5969_o & n5972_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n6004_o = n5969_o & n5976_o;
  assign n6005_o = {1'b1, 1'b1};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n6007_o = n5969_o ? n6005_o : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n6009_o = n5969_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2676:49  */
  assign n6011_o = n5969_o ? n5988_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6012_o = n5822_o ? n5936_o : make_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6013_o = n5822_o ? n5937_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6014_o = n5822_o ? n5938_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6016_o = n5822_o ? n5940_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6017_o = n5822_o ? n5942_o : n5991_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6018_o = n5822_o ? n5944_o : n5994_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6020_o = n5822_o ? n5946_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6021_o = n5822_o ? n5948_o : n5997_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6022_o = n5822_o ? n5950_o : n6000_o;
  assign n6023_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6024_o = n5822_o ? n6023_o : n5975_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6026_o = n5822_o & n5952_o;
  assign n6027_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6028_o = n5822_o ? n6027_o : n5979_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6029_o = n5822_o ? n5953_o : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6031_o = n5822_o ? 2'b00 : n6007_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6033_o = n5822_o ? n5955_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6035_o = n5822_o ? 1'b0 : n6009_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6036_o = n5822_o ? n5957_o : n6011_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2631:41  */
  assign n6037_o = n5822_o ? n5958_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2630:25  */
  assign n6039_o = n2140_o == 4'b0101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:47  */
  assign n6041_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2703:50  */
  assign n6042_o = opcode[11:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2703:63  */
  assign n6044_o = n6042_o == 4'b0001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2706:58  */
  assign n6046_o = opcode[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2706:70  */
  assign n6048_o = n6046_o == 8'b11111111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2709:61  */
  assign n6050_o = opcode[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2709:73  */
  assign n6052_o = n6050_o == 8'b00000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2709:49  */
  assign n6054_o = n6052_o ? n1985_o : 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2709:49  */
  assign n6057_o = n6052_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2709:49  */
  assign n6060_o = n6052_o ? 7'b0010111 : 7'b0010110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2706:49  */
  assign n6061_o = n6048_o ? n1985_o : n6054_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2706:49  */
  assign n6063_o = n6048_o ? 1'b0 : n6057_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2706:49  */
  assign n6064_o = n6048_o ? 1'b1 : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2706:49  */
  assign n6066_o = n6048_o ? 7'b0010111 : n6060_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2717:58  */
  assign n6067_o = opcode[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2717:70  */
  assign n6069_o = n6067_o == 8'b11111111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2720:61  */
  assign n6071_o = opcode[7:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2720:73  */
  assign n6073_o = n6071_o == 8'b00000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2720:49  */
  assign n6075_o = n6073_o ? n1985_o : 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2717:49  */
  assign n6076_o = n6069_o ? n1985_o : n6075_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2717:49  */
  assign n6077_o = n6069_o ? 1'b1 : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2703:41  */
  assign n6078_o = n6044_o ? n6061_o : n6076_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:33  */
  assign n6080_o = n6091_o ? 1'b1 : n1974_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2703:41  */
  assign n6082_o = n6044_o ? n6063_o : 1'b0;
  assign n6083_o = n2121_o[1];
  assign n6084_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n6085_o = n1996_o ? n6083_o : n6084_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2703:41  */
  assign n6086_o = n6044_o ? 1'b1 : n6085_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2703:41  */
  assign n6087_o = n6044_o ? n6064_o : n6077_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2703:41  */
  assign n6089_o = n6044_o ? n6066_o : 7'b0010101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:33  */
  assign n6090_o = n6041_o ? n6078_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:33  */
  assign n6091_o = n6041_o & n6044_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:33  */
  assign n6093_o = n6041_o ? n6082_o : 1'b0;
  assign n6094_o = n2121_o[1];
  assign n6095_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n6096_o = n1996_o ? n6094_o : n6095_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:33  */
  assign n6097_o = n6041_o ? n6086_o : n6096_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:33  */
  assign n6098_o = n6041_o ? n6087_o : n2130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2702:33  */
  assign n6099_o = n6041_o ? n6089_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2699:25  */
  assign n6101_o = n2140_o == 4'b0110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:42  */
  assign n6102_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:45  */
  assign n6103_o = ~n6102_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:33  */
  assign n6108_o = n6103_o ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:33  */
  assign n6111_o = n6103_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:33  */
  assign n6114_o = n6103_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:33  */
  assign n6117_o = n6103_o ? 1'b0 : 1'b1;
  assign n6118_o = {1'b1, 1'b1};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:33  */
  assign n6120_o = n6103_o ? n6118_o : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2731:33  */
  assign n6122_o = n6103_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2730:25  */
  assign n6124_o = n2140_o == 4'b0111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:42  */
  assign n6125_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:54  */
  assign n6127_o = n6125_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:50  */
  assign n6128_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:62  */
  assign n6130_o = n6128_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:56  */
  assign n6132_o = 1'b1 & n6130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:81  */
  assign n6133_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:93  */
  assign n6135_o = n6133_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:111  */
  assign n6136_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:123  */
  assign n6138_o = n6136_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:102  */
  assign n6139_o = n6135_o | n6138_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2746:70  */
  assign n6140_o = n6132_o & n6139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2747:58  */
  assign n6141_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2747:70  */
  assign n6143_o = n6141_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2747:49  */
  assign n6146_o = n6143_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2750:64  */
  assign n6148_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2750:70  */
  assign n6149_o = n6148_o & nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2750:98  */
  assign n6150_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2750:110  */
  assign n6152_o = n6150_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2750:116  */
  assign n6153_o = n6152_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2750:88  */
  assign n6154_o = n6149_o | n6153_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6156_o = n6410_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6158_o = n6194_o ? 7'b1010101 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2755:59  */
  assign n6159_o = ~z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2755:78  */
  assign n6160_o = ~set_v_flag;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2755:64  */
  assign n6161_o = n6159_o & n6160_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2755:49  */
  assign n6164_o = n6161_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2759:75  */
  assign n6165_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2759:87  */
  assign n6167_o = n6165_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2759:93  */
  assign n6168_o = n6167_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2759:65  */
  assign n6169_o = nextpass | n6168_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2759:49  */
  assign n6172_o = n6169_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6174_o = n6140_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6175_o = n6140_o & n6154_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6177_o = n6140_o ? n6146_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6180_o = n6140_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6182_o = n6140_o ? n6172_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6185_o = n6140_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6188_o = n6140_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6191_o = n6140_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6193_o = n6140_o ? n6164_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2745:41  */
  assign n6194_o = n6140_o & n6154_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:45  */
  assign n6195_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:63  */
  assign n6196_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:75  */
  assign n6198_o = n6196_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:53  */
  assign n6199_o = n6195_o & n6198_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:50  */
  assign n6200_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:62  */
  assign n6202_o = n6200_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:53  */
  assign n6206_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:65  */
  assign n6208_o = n6206_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:80  */
  assign n6209_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:92  */
  assign n6211_o = n6209_o == 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:71  */
  assign n6212_o = n6208_o | n6211_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2777:58  */
  assign n6215_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2777:71  */
  assign n6217_o = n6215_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2777:49  */
  assign n6222_o = n6217_o ? 2'b01 : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2777:49  */
  assign n6224_o = n6217_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2777:49  */
  assign n6226_o = n6217_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:58  */
  assign n6227_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:61  */
  assign n6228_o = ~n6227_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2785:66  */
  assign n6229_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2785:79  */
  assign n6231_o = n6229_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2785:57  */
  assign n6234_o = n6231_o ? 2'b00 : 2'b01;
  assign n6238_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6239_o = n6280_o ? 1'b1 : n6238_o;
  assign n6240_o = n1870_o[80];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6241_o = n6284_o ? 1'b1 : n6240_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2792:57  */
  assign n6243_o = decodeopc ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2800:57  */
  assign n6245_o = decodeopc ? 1'b1 : n2113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2800:57  */
  assign n6247_o = decodeopc ? 7'b0011110 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6248_o = n6264_o ? n6234_o : datatype;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:49  */
  assign n6251_o = n6228_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:49  */
  assign n6254_o = n6228_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:49  */
  assign n6255_o = n6228_o ? n2113_o : n6245_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:49  */
  assign n6257_o = n6228_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:49  */
  assign n6259_o = n6228_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:49  */
  assign n6261_o = n6228_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2784:49  */
  assign n6262_o = n6228_o ? n6243_o : n6247_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6263_o = n6212_o ? n6222_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6264_o = n6212_o & n6228_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6266_o = n6212_o ? n6251_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6269_o = n6212_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6271_o = n6212_o ? n6254_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6272_o = n6212_o ? n6255_o : n2113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6275_o = n6212_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6278_o = n6212_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6280_o = n6212_o & n6257_o;
  assign n6281_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6282_o = n6212_o ? 1'b1 : n6281_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6284_o = n6212_o & n6259_o;
  assign n6285_o = {n6226_o, n6224_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6287_o = n6212_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6289_o = n6212_o ? n6261_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6291_o = n6212_o ? n6285_o : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2773:41  */
  assign n6292_o = n6212_o ? n6262_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6293_o = n6202_o ? n1882_o : n6263_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6294_o = n6202_o ? datatype : n6248_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6296_o = n6202_o ? 1'b0 : n6266_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6298_o = n6202_o ? 1'b0 : n6269_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6300_o = n6202_o ? 1'b0 : n6271_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6301_o = n6202_o ? n2113_o : n6272_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6303_o = n6202_o ? 1'b0 : n6275_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6305_o = n6202_o ? 1'b0 : n6278_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6308_o = n6202_o ? 1'b1 : 1'b0;
  assign n6309_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6310_o = n6202_o ? n6309_o : n6239_o;
  assign n6311_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6312_o = n6202_o ? n6311_o : n6282_o;
  assign n6313_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6314_o = n6392_o ? 1'b1 : n6313_o;
  assign n6315_o = n1870_o[80];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6316_o = n6202_o ? n6315_o : n6241_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6318_o = n6202_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6320_o = n6202_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6322_o = n6202_o ? 1'b0 : n6287_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6324_o = n6202_o ? 1'b0 : n6289_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6326_o = n6202_o ? 2'b00 : n6291_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2768:41  */
  assign n6327_o = n6202_o ? n2139_o : n6292_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2810:50  */
  assign n6328_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2810:62  */
  assign n6330_o = n6328_o != 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:52  */
  assign n6331_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:55  */
  assign n6332_o = ~n6331_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:70  */
  assign n6333_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:82  */
  assign n6335_o = n6333_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:60  */
  assign n6336_o = n6332_o & n6335_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:101  */
  assign n6337_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:113  */
  assign n6339_o = n6337_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:131  */
  assign n6340_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:143  */
  assign n6342_o = n6340_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:122  */
  assign n6343_o = n6339_o | n6342_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:90  */
  assign n6344_o = n6336_o & n6343_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:51  */
  assign n6345_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:69  */
  assign n6346_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:81  */
  assign n6348_o = n6346_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:59  */
  assign n6349_o = n6345_o & n6348_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:99  */
  assign n6350_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:111  */
  assign n6352_o = n6350_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:128  */
  assign n6353_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:140  */
  assign n6355_o = n6353_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:119  */
  assign n6356_o = n6352_o | n6355_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2812:88  */
  assign n6357_o = n6349_o & n6356_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2811:151  */
  assign n6358_o = n6344_o | n6357_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2810:69  */
  assign n6359_o = n6330_o & n6358_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2810:41  */
  assign n6363_o = n6359_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2810:41  */
  assign n6366_o = n6359_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2810:41  */
  assign n6369_o = n6359_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2810:41  */
  assign n6371_o = n6359_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6372_o = n6199_o ? n6293_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6373_o = n6199_o ? n6294_o : datatype;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6375_o = n6199_o ? n6296_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6377_o = n6199_o ? n6298_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6379_o = n6199_o ? n6300_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6380_o = n6199_o ? n6301_o : n2113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6381_o = n6199_o ? n6303_o : n6363_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6382_o = n6199_o ? n6305_o : n6366_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6384_o = n6199_o ? 1'b0 : n6369_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6386_o = n6199_o ? n6308_o : 1'b0;
  assign n6387_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6388_o = n6199_o ? n6310_o : n6387_o;
  assign n6389_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6390_o = n6199_o ? n6312_o : n6389_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6392_o = n6199_o & n6202_o;
  assign n6393_o = n1870_o[80];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6394_o = n6199_o ? n6316_o : n6393_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6396_o = n6199_o ? n6318_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6398_o = n6199_o ? 1'b0 : n6371_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6400_o = n6199_o ? n6320_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6402_o = n6199_o ? n6322_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6404_o = n6199_o ? n6324_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6406_o = n6199_o ? n6326_o : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2767:33  */
  assign n6407_o = n6199_o ? n6327_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6408_o = n6127_o ? n6174_o : n6372_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6409_o = n6127_o ? datatype : n6373_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6410_o = n6127_o & n6175_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6412_o = n6127_o ? n6177_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6414_o = n6127_o ? 1'b0 : n6375_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6415_o = n6127_o ? n6180_o : n6377_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6416_o = n6127_o ? n6182_o : n6379_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6417_o = n6127_o ? n2113_o : n6380_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6418_o = n6127_o ? n6185_o : n6381_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6419_o = n6127_o ? n6188_o : n6382_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6421_o = n6127_o ? n6191_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6423_o = n6127_o ? 1'b0 : n6384_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6425_o = n6127_o ? 1'b0 : n6386_o;
  assign n6426_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6427_o = n6127_o ? n6426_o : n6388_o;
  assign n6428_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6429_o = n6127_o ? n6428_o : n6390_o;
  assign n6430_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6431_o = n6127_o ? n6430_o : n6314_o;
  assign n6432_o = n1870_o[80];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6433_o = n6127_o ? n6432_o : n6394_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6435_o = n6127_o ? 1'b0 : n6396_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6437_o = n6127_o ? 1'b0 : n6398_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6439_o = n6127_o ? 1'b0 : n6400_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6441_o = n6127_o ? 1'b0 : n6402_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6442_o = n6127_o ? n6193_o : n6404_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6444_o = n6127_o ? 2'b00 : n6406_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2744:33  */
  assign n6445_o = n6127_o ? n6158_o : n6407_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2743:25  */
  assign n6447_o = n2140_o == 4'b1000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:42  */
  assign n6448_o = opcode[8:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:54  */
  assign n6450_o = n6448_o != 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:45  */
  assign n6451_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:48  */
  assign n6452_o = ~n6451_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:62  */
  assign n6453_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:74  */
  assign n6455_o = n6453_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:53  */
  assign n6456_o = n6452_o | n6455_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:92  */
  assign n6457_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:104  */
  assign n6459_o = n6457_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:122  */
  assign n6460_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:134  */
  assign n6462_o = n6460_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:113  */
  assign n6463_o = n6459_o | n6462_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:81  */
  assign n6464_o = n6456_o & n6463_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2825:43  */
  assign n6465_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2825:62  */
  assign n6466_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2825:74  */
  assign n6468_o = n6466_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2825:91  */
  assign n6469_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2825:103  */
  assign n6471_o = n6469_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2825:82  */
  assign n6472_o = n6468_o | n6471_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2825:51  */
  assign n6473_o = n6465_o & n6472_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2824:142  */
  assign n6474_o = n6464_o | n6473_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:65  */
  assign n6475_o = n6450_o & n6474_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2828:50  */
  assign n6477_o = opcode[14];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2828:54  */
  assign n6478_o = ~n6477_o;
  assign n6480_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6481_o = n6555_o ? 1'b1 : n6480_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:50  */
  assign n6482_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:62  */
  assign n6484_o = n6482_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2832:58  */
  assign n6485_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2832:61  */
  assign n6486_o = ~n6485_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6488_o = n6530_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2837:58  */
  assign n6490_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2837:49  */
  assign n6493_o = n6490_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2841:49  */
  assign n6497_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2841:49  */
  assign n6500_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2846:58  */
  assign n6501_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2846:76  */
  assign n6502_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2846:88  */
  assign n6504_o = n6502_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2846:66  */
  assign n6505_o = n6501_o & n6504_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2846:49  */
  assign n6508_o = n6505_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2846:49  */
  assign n6511_o = n6505_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6512_o = n6484_o & n6486_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6514_o = n6484_o ? n6493_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6517_o = n6484_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6519_o = n6484_o ? n6497_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6521_o = n6484_o ? n6500_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6523_o = n6484_o ? 1'b0 : n6508_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6525_o = n6484_o ? 1'b0 : n6511_o;
  assign n6526_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6527_o = n6553_o ? 1'b1 : n6526_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2831:41  */
  assign n6529_o = n6484_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6530_o = n6475_o & n6512_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6532_o = n6475_o ? n6514_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6534_o = n6475_o ? n6517_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6536_o = n6475_o ? n6519_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6538_o = n6475_o ? n6521_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6541_o = n6475_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6544_o = n6475_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6547_o = n6475_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6549_o = n6475_o ? n6523_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6551_o = n6475_o ? n6525_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6553_o = n6475_o & n6484_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6555_o = n6475_o & n6478_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6557_o = n6475_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2823:33  */
  assign n6559_o = n6475_o ? n6529_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2822:25  */
  assign n6561_o = n2140_o == 4'b1001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2822:36  */
  assign n6563_o = n2140_o == 4'b1101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2822:36  */
  assign n6564_o = n6561_o | n6563_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2858:25  */
  assign n6566_o = n2140_o == 4'b1010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:42  */
  assign n6567_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:54  */
  assign n6569_o = n6567_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:50  */
  assign n6570_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:62  */
  assign n6572_o = n6570_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:80  */
  assign n6573_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:92  */
  assign n6575_o = n6573_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:71  */
  assign n6576_o = n6572_o | n6575_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2866:58  */
  assign n6577_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2866:61  */
  assign n6578_o = ~n6577_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6581_o = n6745_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2866:49  */
  assign n6583_o = n6578_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2873:66  */
  assign n6585_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2873:57  */
  assign n6588_o = n6585_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2871:49  */
  assign n6590_o = setexecopc ? n6588_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2871:49  */
  assign n6593_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2871:49  */
  assign n6596_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2871:49  */
  assign n6599_o = setexecopc ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6601_o = n6576_o & n6578_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6603_o = n6576_o ? n6590_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6605_o = n6576_o ? n6593_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6607_o = n6576_o ? n6596_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6609_o = n6576_o ? n6599_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6612_o = n6576_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6615_o = n6576_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6618_o = n6576_o ? 1'b1 : 1'b0;
  assign n6619_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6620_o = n6576_o ? 1'b1 : n6619_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6622_o = n6576_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2864:41  */
  assign n6624_o = n6576_o ? n6583_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:50  */
  assign n6625_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:58  */
  assign n6626_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:70  */
  assign n6628_o = n6626_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2890:74  */
  assign n6630_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2890:86  */
  assign n6632_o = n6630_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6634_o = n6734_o ? 1'b1 : n2127_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6638_o = n6724_o ? 2'b10 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6639_o = n6729_o ? 1'b1 : n1966_o;
  assign n6640_o = n2121_o[0];
  assign n6641_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n6642_o = n1996_o ? n6640_o : n6641_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2889:57  */
  assign n6643_o = decodeopc ? 1'b1 : n6642_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2889:57  */
  assign n6644_o = decodeopc & n6632_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6646_o = n6744_o ? 7'b0100010 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:66  */
  assign n6649_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:78  */
  assign n6651_o = n6649_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:95  */
  assign n6652_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:107  */
  assign n6654_o = n6652_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:86  */
  assign n6655_o = n6651_o | n6654_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:57  */
  assign n6659_o = n6655_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:57  */
  assign n6662_o = n6655_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:57  */
  assign n6665_o = n6655_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:57  */
  assign n6668_o = n6655_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2901:57  */
  assign n6670_o = n6655_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6671_o = n6628_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6673_o = n6628_o ? 1'b0 : n6659_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6675_o = n6628_o ? 1'b0 : n6662_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6677_o = n6628_o ? 1'b1 : n6665_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6679_o = n6628_o ? 1'b0 : n6668_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6680_o = n6628_o & decodeopc;
  assign n6681_o = n2121_o[0];
  assign n6682_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n6683_o = n1996_o ? n6681_o : n6682_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6684_o = n6628_o ? n6643_o : n6683_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6685_o = n6628_o & n6644_o;
  assign n6686_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6687_o = n6628_o ? 1'b1 : n6686_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6689_o = n6628_o ? 1'b0 : n6670_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6691_o = n6628_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6693_o = n6628_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2886:49  */
  assign n6694_o = n6628_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:58  */
  assign n6695_o = opcode[8:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:70  */
  assign n6697_o = n6695_o != 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2912:59  */
  assign n6698_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2912:71  */
  assign n6700_o = n6698_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2912:89  */
  assign n6701_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2912:101  */
  assign n6703_o = n6701_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2912:80  */
  assign n6704_o = n6700_o | n6703_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:81  */
  assign n6705_o = n6697_o & n6704_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:49  */
  assign n6710_o = n6705_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:49  */
  assign n6713_o = n6705_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:49  */
  assign n6716_o = n6705_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:49  */
  assign n6719_o = n6705_o ? 1'b1 : 1'b0;
  assign n6720_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:49  */
  assign n6721_o = n6705_o ? 1'b1 : n6720_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2911:49  */
  assign n6723_o = n6705_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6724_o = n6625_o & n6671_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6725_o = n6625_o ? n6673_o : n6710_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6726_o = n6625_o ? n6675_o : n6713_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6727_o = n6625_o ? n6677_o : n6716_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6728_o = n6625_o ? n6679_o : n6719_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6729_o = n6625_o & n6680_o;
  assign n6730_o = n2121_o[0];
  assign n6731_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n6732_o = n1996_o ? n6730_o : n6731_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6733_o = n6625_o ? n6684_o : n6732_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6734_o = n6625_o & n6685_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6735_o = n6625_o ? n6687_o : n6721_o;
  assign n6736_o = {n6691_o, n6689_o};
  assign n6737_o = n6736_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6739_o = n6625_o ? n6737_o : 1'b0;
  assign n6740_o = n6736_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6741_o = n6625_o ? n6740_o : n6723_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6743_o = n6625_o ? n6693_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2885:41  */
  assign n6744_o = n6625_o & n6694_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6745_o = n6569_o & n6601_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6746_o = n6569_o ? n1985_o : n6638_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6748_o = n6569_o ? n6603_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6750_o = n6569_o ? n6605_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6752_o = n6569_o ? n6607_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6754_o = n6569_o ? n6609_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6755_o = n6569_o ? n6612_o : n6725_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6756_o = n6569_o ? n6615_o : n6726_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6757_o = n6569_o ? n6618_o : n6727_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6759_o = n6569_o ? 1'b0 : n6728_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6760_o = n6569_o ? n1966_o : n6639_o;
  assign n6761_o = n2121_o[0];
  assign n6762_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n6763_o = n1996_o ? n6761_o : n6762_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6764_o = n6569_o ? n6763_o : n6733_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6765_o = n6569_o ? n2127_o : n6634_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6766_o = n6569_o ? n6620_o : n6735_o;
  assign n6767_o = {n6741_o, n6739_o};
  assign n6768_o = n6767_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6770_o = n6569_o ? 1'b0 : n6768_o;
  assign n6771_o = n6767_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6772_o = n6569_o ? n6622_o : n6771_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6774_o = n6569_o ? n6624_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6776_o = n6569_o ? 1'b0 : n6743_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2863:33  */
  assign n6777_o = n6569_o ? n2139_o : n6646_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2862:25  */
  assign n6779_o = n2140_o == 4'b1011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:42  */
  assign n6780_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:54  */
  assign n6782_o = n6780_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:50  */
  assign n6783_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:62  */
  assign n6785_o = n6783_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:56  */
  assign n6787_o = 1'b1 & n6785_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:81  */
  assign n6788_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:93  */
  assign n6790_o = n6788_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:111  */
  assign n6791_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:123  */
  assign n6793_o = n6791_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:102  */
  assign n6794_o = n6790_o | n6793_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2928:70  */
  assign n6795_o = n6787_o & n6794_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2929:58  */
  assign n6796_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2929:70  */
  assign n6798_o = n6796_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2929:49  */
  assign n6801_o = n6798_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:64  */
  assign n6803_o = micro_state == 7'b0000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:70  */
  assign n6804_o = n6803_o & nextpass;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:98  */
  assign n6805_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:110  */
  assign n6807_o = n6805_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:116  */
  assign n6808_o = n6807_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:88  */
  assign n6809_o = n6804_o | n6808_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:49  */
  assign n6813_o = n6809_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2932:49  */
  assign n6815_o = n6809_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2945:77  */
  assign n6817_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2945:89  */
  assign n6819_o = n6817_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2945:95  */
  assign n6820_o = n6819_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2945:67  */
  assign n6821_o = nextpass | n6820_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2945:49  */
  assign n6824_o = n6821_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2949:49  */
  assign n6827_o = setexecopc ? 2'b10 : 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6829_o = n6795_o ? n6827_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6831_o = n6795_o ? n6801_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6834_o = n6795_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6836_o = n6795_o ? n6824_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6839_o = n6795_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6842_o = n6795_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6845_o = n6795_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6847_o = n6795_o ? n6813_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6849_o = n6795_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2927:41  */
  assign n6851_o = n6795_o ? n6815_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:45  */
  assign n6852_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:63  */
  assign n6853_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:75  */
  assign n6855_o = n6853_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:53  */
  assign n6856_o = n6852_o & n6855_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:50  */
  assign n6857_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:62  */
  assign n6859_o = n6857_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:58  */
  assign n6862_o = opcode[7:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:70  */
  assign n6864_o = n6862_o == 4'b0100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:87  */
  assign n6865_o = opcode[7:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:99  */
  assign n6867_o = n6865_o == 5'b10001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:78  */
  assign n6868_o = n6864_o | n6867_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2967:66  */
  assign n6872_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2967:84  */
  assign n6873_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2967:74  */
  assign n6874_o = n6872_o & n6873_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2967:57  */
  assign n6877_o = n6874_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2967:57  */
  assign n6880_o = n6874_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6882_o = n6888_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2971:57  */
  assign n6885_o = decodeopc ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6887_o = n6868_o ? 2'b10 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6888_o = n6868_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6890_o = n6868_o ? n6877_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6892_o = n6868_o ? n6880_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6894_o = n6868_o ? n6885_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6897_o = n6868_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6900_o = n6868_o ? 1'b0 : 1'b1;
  assign n6901_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6902_o = n6868_o ? 1'b1 : n6901_o;
  assign n6903_o = n1870_o[61];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6904_o = n6868_o ? 1'b1 : n6903_o;
  assign n6905_o = n1870_o[85];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2962:49  */
  assign n6906_o = n6868_o ? 1'b1 : n6905_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6907_o = n6859_o ? n1882_o : n6887_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6908_o = n6859_o ? n1985_o : n6882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6910_o = n6859_o ? 1'b0 : n6890_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6912_o = n6859_o ? 1'b0 : n6892_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6914_o = n6859_o ? 1'b0 : n6894_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6916_o = n6859_o ? 1'b0 : n6897_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6918_o = n6859_o ? 1'b0 : n6900_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6921_o = n6859_o ? 1'b1 : 1'b0;
  assign n6922_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6923_o = n6859_o ? n6922_o : n6902_o;
  assign n6924_o = n1870_o[61];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6925_o = n6859_o ? n6924_o : n6904_o;
  assign n6926_o = n1870_o[85];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6927_o = n6859_o ? n6926_o : n6906_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6929_o = n6859_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2957:41  */
  assign n6931_o = n6859_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2982:50  */
  assign n6932_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2982:62  */
  assign n6934_o = n6932_o != 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:52  */
  assign n6935_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:55  */
  assign n6936_o = ~n6935_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:70  */
  assign n6937_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:82  */
  assign n6939_o = n6937_o != 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:60  */
  assign n6940_o = n6936_o & n6939_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:101  */
  assign n6941_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:113  */
  assign n6943_o = n6941_o != 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:131  */
  assign n6944_o = opcode[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:143  */
  assign n6946_o = n6944_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:122  */
  assign n6947_o = n6943_o | n6946_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:90  */
  assign n6948_o = n6940_o & n6947_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:51  */
  assign n6949_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:69  */
  assign n6950_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:81  */
  assign n6952_o = n6950_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:59  */
  assign n6953_o = n6949_o & n6952_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:99  */
  assign n6954_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:111  */
  assign n6956_o = n6954_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:128  */
  assign n6957_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:140  */
  assign n6959_o = n6957_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:119  */
  assign n6960_o = n6956_o | n6959_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2984:88  */
  assign n6961_o = n6953_o & n6960_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2983:151  */
  assign n6962_o = n6948_o | n6961_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2982:69  */
  assign n6963_o = n6934_o & n6962_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2982:41  */
  assign n6967_o = n6963_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2982:41  */
  assign n6970_o = n6963_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2982:41  */
  assign n6973_o = n6963_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2982:41  */
  assign n6975_o = n6963_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6976_o = n6856_o ? n6907_o : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6977_o = n6856_o ? n6908_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6979_o = n6856_o ? n6910_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6981_o = n6856_o ? n6912_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6983_o = n6856_o ? n6914_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6984_o = n6856_o ? n6916_o : n6967_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6985_o = n6856_o ? n6918_o : n6970_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6987_o = n6856_o ? 1'b0 : n6973_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6989_o = n6856_o ? n6921_o : 1'b0;
  assign n6990_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6991_o = n6856_o ? n6923_o : n6990_o;
  assign n6992_o = n1870_o[61];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6993_o = n6856_o ? n6925_o : n6992_o;
  assign n6994_o = n1870_o[85];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6995_o = n6856_o ? n6927_o : n6994_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6997_o = n6856_o ? n6929_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n6999_o = n6856_o ? 1'b0 : n6975_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2956:33  */
  assign n7001_o = n6856_o ? n6931_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7002_o = n6782_o ? n6829_o : n6976_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7003_o = n6782_o ? n1985_o : n6977_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7005_o = n6782_o ? n6831_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7007_o = n6782_o ? 1'b0 : n6979_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7009_o = n6782_o ? n6834_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7011_o = n6782_o ? 1'b0 : n6981_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7012_o = n6782_o ? n6836_o : n6983_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7013_o = n6782_o ? n6839_o : n6984_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7014_o = n6782_o ? n6842_o : n6985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7016_o = n6782_o ? n6845_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7018_o = n6782_o ? 1'b0 : n6987_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7020_o = n6782_o ? 1'b0 : n6989_o;
  assign n7021_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7022_o = n6782_o ? n7021_o : n6991_o;
  assign n7023_o = n1870_o[61];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7024_o = n6782_o ? n7023_o : n6993_o;
  assign n7025_o = n1870_o[85];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7026_o = n6782_o ? n7025_o : n6995_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7028_o = n6782_o ? 1'b0 : n6997_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7030_o = n6782_o ? 1'b0 : n6999_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7032_o = n6782_o ? 1'b0 : n7001_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7034_o = n6782_o ? n6847_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7036_o = n6782_o ? n6849_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2926:33  */
  assign n7038_o = n6782_o ? n6851_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2925:25  */
  assign n7040_o = n2140_o == 4'b1100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:42  */
  assign n7041_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:54  */
  assign n7043_o = n7041_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:50  */
  assign n7044_o = opcode[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:54  */
  assign n7045_o = ~n7044_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:54  */
  assign n7046_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:66  */
  assign n7048_o = n7046_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:84  */
  assign n7049_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:96  */
  assign n7051_o = n7049_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:113  */
  assign n7052_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:125  */
  assign n7054_o = n7052_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:104  */
  assign n7055_o = n7051_o | n7054_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:73  */
  assign n7056_o = n7048_o & n7055_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3005:79  */
  assign n7058_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7061_o = n7346_o ? 2'b01 : n1882_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:44  */
  assign n7064_o = n7056_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7065_o = n7363_o ? n7058_o : n1861_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:44  */
  assign n7068_o = n7056_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:44  */
  assign n7071_o = n7056_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:44  */
  assign n7074_o = n7056_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:44  */
  assign n7076_o = n7056_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2997:44  */
  assign n7078_o = n7056_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:70  */
  assign n7079_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:73  */
  assign n7080_o = ~n7079_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:78  */
  assign n7082_o = n7080_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:63  */
  assign n7084_o = 1'b0 | n7082_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:60  */
  assign n7085_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:73  */
  assign n7087_o = n7085_o == 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:88  */
  assign n7088_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:101  */
  assign n7090_o = n7088_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:79  */
  assign n7091_o = n7087_o | n7090_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:117  */
  assign n7092_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:130  */
  assign n7094_o = n7092_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:108  */
  assign n7095_o = n7091_o | n7094_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:59  */
  assign n7096_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:71  */
  assign n7098_o = n7096_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:87  */
  assign n7099_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:99  */
  assign n7101_o = n7099_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:78  */
  assign n7102_o = n7098_o | n7101_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:115  */
  assign n7103_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:127  */
  assign n7105_o = n7103_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:106  */
  assign n7106_o = n7102_o | n7105_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:144  */
  assign n7107_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:156  */
  assign n7109_o = n7107_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:173  */
  assign n7110_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:185  */
  assign n7112_o = n7110_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:163  */
  assign n7113_o = n7109_o & n7112_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:134  */
  assign n7114_o = n7106_o | n7113_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3014:138  */
  assign n7115_o = n7095_o & n7114_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:94  */
  assign n7116_o = n7084_o | n7115_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:60  */
  assign n7117_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:73  */
  assign n7119_o = n7117_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:88  */
  assign n7120_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:101  */
  assign n7122_o = n7120_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:79  */
  assign n7123_o = n7119_o | n7122_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:117  */
  assign n7124_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:130  */
  assign n7126_o = n7124_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:108  */
  assign n7127_o = n7123_o | n7126_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:59  */
  assign n7128_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:71  */
  assign n7130_o = n7128_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:87  */
  assign n7131_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:99  */
  assign n7133_o = n7131_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:78  */
  assign n7134_o = n7130_o | n7133_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:115  */
  assign n7135_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:127  */
  assign n7137_o = n7135_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:106  */
  assign n7138_o = n7134_o | n7137_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:143  */
  assign n7139_o = opcode[5:2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:155  */
  assign n7141_o = n7139_o == 4'b1111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3017:134  */
  assign n7142_o = n7138_o | n7141_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3016:138  */
  assign n7143_o = n7127_o & n7142_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3015:195  */
  assign n7144_o = n7116_o | n7143_o;
  assign n7147_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3021:57  */
  assign n7148_o = decodeopc ? 1'b1 : n7147_o;
  assign n7149_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3021:57  */
  assign n7150_o = decodeopc ? 1'b1 : n7149_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3021:57  */
  assign n7152_o = decodeopc ? 7'b0000001 : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3028:66  */
  assign n7154_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3028:84  */
  assign n7155_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3028:87  */
  assign n7156_o = ~n7155_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3028:75  */
  assign n7157_o = n7154_o | n7156_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3028:57  */
  assign n7160_o = n7157_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3031:66  */
  assign n7161_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3031:79  */
  assign n7163_o = n7161_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3031:57  */
  assign n7166_o = n7163_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:66  */
  assign n7167_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:79  */
  assign n7169_o = n7167_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:95  */
  assign n7170_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:108  */
  assign n7172_o = n7170_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:86  */
  assign n7173_o = n7169_o | n7172_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:124  */
  assign n7174_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:137  */
  assign n7176_o = n7174_o == 3'b110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:115  */
  assign n7177_o = n7173_o | n7176_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:153  */
  assign n7178_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:166  */
  assign n7180_o = n7178_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:144  */
  assign n7181_o = n7177_o | n7180_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3034:57  */
  assign n7184_o = n7181_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:66  */
  assign n7185_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:79  */
  assign n7187_o = n7185_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:95  */
  assign n7188_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:108  */
  assign n7190_o = n7188_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:86  */
  assign n7191_o = n7187_o | n7190_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:124  */
  assign n7192_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:137  */
  assign n7194_o = n7192_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:115  */
  assign n7195_o = n7191_o | n7194_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3038:57  */
  assign n7198_o = n7195_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:66  */
  assign n7199_o = opcode[4:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:78  */
  assign n7201_o = n7199_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3042:74  */
  assign n7202_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3042:87  */
  assign n7204_o = n7202_o != 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7206_o = n7226_o ? 1'b1 : n7198_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3045:72  */
  assign n7207_o = exec[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7210_o = n7219_o ? 2'b01 : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3045:65  */
  assign n7213_o = n7207_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3045:65  */
  assign n7216_o = n7207_o ? 1'b1 : 1'b0;
  assign n7217_o = n1870_o[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7218_o = n7225_o ? 1'b1 : n7217_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7219_o = n7201_o & n7207_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7221_o = n7201_o ? n7213_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7223_o = n7201_o ? n7216_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7225_o = n7201_o & n7207_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3041:57  */
  assign n7226_o = n7201_o & n7204_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3052:63  */
  assign n7227_o = set[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3052:57  */
  assign n7229_o = n7227_o ? 2'b01 : n7210_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3055:64  */
  assign n7230_o = exec[62];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3055:57  */
  assign n7234_o = n7230_o ? 2'b01 : n7229_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3055:57  */
  assign n7236_o = n7230_o ? 1'b1 : n7221_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3055:57  */
  assign n7238_o = n7230_o ? 1'b1 : n7223_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3055:57  */
  assign n7239_o = n7230_o ? 1'b1 : n7218_o;
  assign n7240_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3055:57  */
  assign n7241_o = n7230_o ? 1'b1 : n7240_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3055:57  */
  assign n7243_o = n7230_o ? 7'b1010000 : n7152_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3064:74  */
  assign n7244_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3064:87  */
  assign n7246_o = n7244_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3064:65  */
  assign n7249_o = n7246_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3064:65  */
  assign n7252_o = n7246_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:74  */
  assign n7253_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:87  */
  assign n7255_o = n7253_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:103  */
  assign n7256_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:116  */
  assign n7258_o = n7256_o == 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:94  */
  assign n7259_o = n7255_o | n7258_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:132  */
  assign n7260_o = opcode[10:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:145  */
  assign n7262_o = n7260_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3069:123  */
  assign n7263_o = n7259_o | n7262_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3063:57  */
  assign n7265_o = n7270_o ? 1'b1 : n7238_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3063:57  */
  assign n7267_o = setexecopc ? n7249_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3063:57  */
  assign n7269_o = setexecopc ? n7252_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3063:57  */
  assign n7270_o = setexecopc & n7263_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7271_o = n7144_o ? n1985_o : n7234_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7273_o = n7144_o ? 1'b0 : n7184_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7276_o = n7144_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7278_o = n7144_o ? 1'b0 : n7267_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7280_o = n7144_o ? 1'b0 : n7269_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7282_o = n7144_o ? 1'b0 : n7236_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7284_o = n7144_o ? 1'b0 : n7265_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7287_o = n7144_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7290_o = n7144_o ? 1'b1 : 1'b0;
  assign n7291_o = n1870_o[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7292_o = n7144_o ? n7291_o : n7239_o;
  assign n7293_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7294_o = n7144_o ? n7293_o : n7148_o;
  assign n7295_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7296_o = n7144_o ? n7295_o : n7241_o;
  assign n7297_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7298_o = n7144_o ? n7297_o : n7150_o;
  assign n7299_o = {n7160_o, 1'b1};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7301_o = n7144_o ? 1'b0 : n7166_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7303_o = n7144_o ? 1'b0 : n7206_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7305_o = n7144_o ? 2'b00 : n7299_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3013:49  */
  assign n7306_o = n7144_o ? n2139_o : n7243_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7307_o = n7045_o & n7056_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7308_o = n7045_o ? n1985_o : n7271_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7309_o = n7045_o ? n7064_o : n7273_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7311_o = n7045_o ? 1'b0 : n7276_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7313_o = n7045_o ? 1'b0 : n7278_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7315_o = n7045_o ? 1'b0 : n7280_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7317_o = n7045_o ? 1'b0 : n7282_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7319_o = n7045_o ? 1'b0 : n7284_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7320_o = n7045_o & n7056_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7321_o = n7045_o ? n7068_o : n7287_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7322_o = n7045_o ? n7071_o : n7290_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7324_o = n7045_o ? n7074_o : 1'b0;
  assign n7325_o = n1870_o[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7326_o = n7045_o ? n7325_o : n7292_o;
  assign n7327_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7328_o = n7045_o ? n7327_o : n7294_o;
  assign n7329_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7330_o = n7045_o ? n7329_o : n7296_o;
  assign n7331_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7332_o = n7045_o ? n7331_o : n7298_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7333_o = n7045_o ? n7076_o : n7301_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7335_o = n7045_o ? 1'b0 : n7303_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7337_o = n7045_o ? 2'b00 : n7305_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7339_o = n7045_o ? n7078_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2996:41  */
  assign n7340_o = n7045_o ? n2139_o : n7306_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7346_o = n7043_o & n7307_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7347_o = n7043_o ? n7308_o : n1985_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7350_o = n7043_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7352_o = n7043_o ? n7309_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7354_o = n7043_o ? n7311_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7356_o = n7043_o ? n7313_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7358_o = n7043_o ? n7315_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7360_o = n7043_o ? n7317_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7362_o = n7043_o ? n7319_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7363_o = n7043_o & n7320_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7365_o = n7043_o ? n7321_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7367_o = n7043_o ? n7322_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7369_o = n7043_o ? n7324_o : 1'b0;
  assign n7370_o = n1870_o[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7371_o = n7043_o ? n7326_o : n7370_o;
  assign n7372_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7373_o = n7043_o ? n7328_o : n7372_o;
  assign n7374_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7375_o = n7043_o ? n7330_o : n7374_o;
  assign n7376_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7377_o = n7043_o ? n7332_o : n7376_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7379_o = n7043_o ? n7333_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7380_o = n7043_o ? n7335_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7382_o = n7043_o ? n7337_o : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7383_o = n7043_o ? n7339_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2995:33  */
  assign n7384_o = n7043_o ? n7340_o : n2139_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:2994:25  */
  assign n7386_o = n2140_o == 4'b1110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3104:39  */
  assign n7387_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3104:57  */
  assign n7388_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3104:69  */
  assign n7390_o = n7388_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3104:47  */
  assign n7391_o = n7387_o & n7390_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:50  */
  assign n7392_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:62  */
  assign n7394_o = n7392_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:79  */
  assign n7395_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:91  */
  assign n7397_o = n7395_o != 3'b011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:69  */
  assign n7398_o = n7394_o & n7397_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3106:51  */
  assign n7399_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3106:63  */
  assign n7401_o = n7399_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3106:80  */
  assign n7402_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3106:92  */
  assign n7404_o = n7402_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3106:71  */
  assign n7405_o = n7401_o | n7404_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:99  */
  assign n7406_o = n7398_o & n7405_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3107:58  */
  assign n7407_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3107:71  */
  assign n7409_o = n7407_o != 3'b000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3109:74  */
  assign n7410_o = opcode[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3109:77  */
  assign n7411_o = ~n7410_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3109:92  */
  assign n7412_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3109:104  */
  assign n7414_o = n7412_o != 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3109:82  */
  assign n7415_o = n7411_o & n7414_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3109:65  */
  assign n7418_o = n7415_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3109:65  */
  assign n7421_o = n7415_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3108:57  */
  assign n7423_o = svmode ? n7418_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3108:57  */
  assign n7426_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3108:57  */
  assign n7428_o = svmode ? n7421_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3123:57  */
  assign n7431_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3123:57  */
  assign n7434_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3107:49  */
  assign n7436_o = n7409_o ? n7423_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3107:49  */
  assign n7437_o = n7409_o ? n7426_o : n7431_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3107:49  */
  assign n7438_o = n7409_o ? n7428_o : n7434_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:41  */
  assign n7440_o = n7406_o ? n7436_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:41  */
  assign n7442_o = n7406_o ? n7437_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3105:41  */
  assign n7444_o = n7406_o ? n7438_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3135:42  */
  assign n7445_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3135:60  */
  assign n7446_o = opcode[8:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3135:72  */
  assign n7448_o = n7446_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3135:50  */
  assign n7449_o = n7445_o & n7448_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:50  */
  assign n7450_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:62  */
  assign n7452_o = n7450_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:79  */
  assign n7453_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:91  */
  assign n7455_o = n7453_o != 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:69  */
  assign n7456_o = n7452_o & n7455_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3137:51  */
  assign n7457_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3137:63  */
  assign n7459_o = n7457_o != 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3137:81  */
  assign n7460_o = opcode[2:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3137:93  */
  assign n7462_o = n7460_o != 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3138:50  */
  assign n7463_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3138:62  */
  assign n7465_o = n7463_o != 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3137:100  */
  assign n7466_o = n7462_o & n7465_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3137:71  */
  assign n7467_o = n7459_o | n7466_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:99  */
  assign n7468_o = n7456_o & n7467_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3139:58  */
  assign n7469_o = opcode[5:1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3139:70  */
  assign n7471_o = n7469_o != 5'b11110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:66  */
  assign n7472_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:79  */
  assign n7474_o = n7472_o == 3'b001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:95  */
  assign n7475_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:108  */
  assign n7477_o = n7475_o == 3'b010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:86  */
  assign n7478_o = n7474_o | n7477_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3142:82  */
  assign n7479_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3142:94  */
  assign n7481_o = n7479_o == 3'b101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3142:73  */
  assign n7484_o = n7481_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3142:73  */
  assign n7487_o = n7481_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3141:65  */
  assign n7489_o = svmode ? n7484_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3141:65  */
  assign n7492_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3141:65  */
  assign n7494_o = svmode ? n7487_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3155:65  */
  assign n7497_o = svmode ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3155:65  */
  assign n7500_o = svmode ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:57  */
  assign n7502_o = n7478_o ? n7489_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:57  */
  assign n7503_o = n7478_o ? n7492_o : n7497_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3140:57  */
  assign n7504_o = n7478_o ? n7494_o : n7500_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3139:49  */
  assign n7506_o = n7471_o ? n7502_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3139:49  */
  assign n7508_o = n7471_o ? n7503_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3139:49  */
  assign n7510_o = n7471_o ? n7504_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:41  */
  assign n7512_o = n7468_o ? n7506_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:41  */
  assign n7514_o = n7468_o ? n7508_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3136:41  */
  assign n7516_o = n7468_o ? n7510_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3135:33  */
  assign n7518_o = n7449_o ? n7512_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3135:33  */
  assign n7520_o = n7449_o ? n7514_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3135:33  */
  assign n7522_o = n7449_o ? n7516_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3104:33  */
  assign n7523_o = n7391_o ? n7440_o : n7518_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3104:33  */
  assign n7524_o = n7391_o ? n7442_o : n7520_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3104:33  */
  assign n7525_o = n7391_o ? n7444_o : n7522_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3103:25  */
  assign n7527_o = n2140_o == 4'b1111;
  assign n7528_o = {n7527_o, n7386_o, n7040_o, n6779_o, n6566_o, n6564_o, n6447_o, n6124_o, n6101_o, n6039_o, n5819_o, n3310_o, n3096_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7529_o = make_berr;
      13'b0100000000000: n7529_o = make_berr;
      13'b0010000000000: n7529_o = make_berr;
      13'b0001000000000: n7529_o = make_berr;
      13'b0000100000000: n7529_o = make_berr;
      13'b0000010000000: n7529_o = make_berr;
      13'b0000001000000: n7529_o = make_berr;
      13'b0000000100000: n7529_o = make_berr;
      13'b0000000010000: n7529_o = make_berr;
      13'b0000000001000: n7529_o = n6012_o;
      13'b0000000000100: n7529_o = n5707_o;
      13'b0000000000010: n7529_o = make_berr;
      13'b0000000000001: n7529_o = make_berr;
      default: n7529_o = make_berr;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7531_o = n1882_o;
      13'b0100000000000: n7531_o = n7061_o;
      13'b0010000000000: n7531_o = n7002_o;
      13'b0001000000000: n7531_o = n6581_o;
      13'b0000100000000: n7531_o = n1882_o;
      13'b0000010000000: n7531_o = n6488_o;
      13'b0000001000000: n7531_o = n6408_o;
      13'b0000000100000: n7531_o = n6108_o;
      13'b0000000010000: n7531_o = 2'b10;
      13'b0000000001000: n7531_o = n6013_o;
      13'b0000000000100: n7531_o = n5708_o;
      13'b0000000000010: n7531_o = n3269_o;
      13'b0000000000001: n7531_o = n3035_o;
      default: n7531_o = n1882_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7532_o = datatype;
      13'b0100000000000: n7532_o = datatype;
      13'b0010000000000: n7532_o = datatype;
      13'b0001000000000: n7532_o = datatype;
      13'b0000100000000: n7532_o = datatype;
      13'b0000010000000: n7532_o = datatype;
      13'b0000001000000: n7532_o = n6409_o;
      13'b0000000100000: n7532_o = datatype;
      13'b0000000010000: n7532_o = datatype;
      13'b0000000001000: n7532_o = datatype;
      13'b0000000000100: n7532_o = datatype;
      13'b0000000000010: n7532_o = datatype;
      13'b0000000000001: n7532_o = datatype;
      default: n7532_o = datatype;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7533_o = n1985_o;
      13'b0100000000000: n7533_o = n7347_o;
      13'b0010000000000: n7533_o = n7003_o;
      13'b0001000000000: n7533_o = n6746_o;
      13'b0000100000000: n7533_o = n1985_o;
      13'b0000010000000: n7533_o = n1985_o;
      13'b0000001000000: n7533_o = n6156_o;
      13'b0000000100000: n7533_o = n1985_o;
      13'b0000000010000: n7533_o = n6090_o;
      13'b0000000001000: n7533_o = n6014_o;
      13'b0000000000100: n7533_o = n5709_o;
      13'b0000000000010: n7533_o = n3259_o;
      13'b0000000000001: n7533_o = n3036_o;
      default: n7533_o = n1985_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7534_o = n2107_o;
      13'b0100000000000: n7534_o = n2107_o;
      13'b0010000000000: n7534_o = n2107_o;
      13'b0001000000000: n7534_o = n2107_o;
      13'b0000100000000: n7534_o = n2107_o;
      13'b0000010000000: n7534_o = n2107_o;
      13'b0000001000000: n7534_o = n2107_o;
      13'b0000000100000: n7534_o = n2107_o;
      13'b0000000010000: n7534_o = n2107_o;
      13'b0000000001000: n7534_o = n2107_o;
      13'b0000000000100: n7534_o = n5710_o;
      13'b0000000000010: n7534_o = n2107_o;
      13'b0000000000001: n7534_o = n2107_o;
      default: n7534_o = n2107_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7536_o = 1'b0;
      13'b0100000000000: n7536_o = 1'b0;
      13'b0010000000000: n7536_o = n7005_o;
      13'b0001000000000: n7536_o = 1'b0;
      13'b0000100000000: n7536_o = 1'b0;
      13'b0000010000000: n7536_o = 1'b0;
      13'b0000001000000: n7536_o = n6412_o;
      13'b0000000100000: n7536_o = 1'b0;
      13'b0000000010000: n7536_o = 1'b0;
      13'b0000000001000: n7536_o = 1'b0;
      13'b0000000000100: n7536_o = 1'b0;
      13'b0000000000010: n7536_o = 1'b0;
      13'b0000000000001: n7536_o = 1'b0;
      default: n7536_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7538_o = n2110_o;
      13'b0100000000000: n7538_o = n2110_o;
      13'b0010000000000: n7538_o = n2110_o;
      13'b0001000000000: n7538_o = n2110_o;
      13'b0000100000000: n7538_o = n2110_o;
      13'b0000010000000: n7538_o = n2110_o;
      13'b0000001000000: n7538_o = n2110_o;
      13'b0000000100000: n7538_o = n2110_o;
      13'b0000000010000: n7538_o = n2110_o;
      13'b0000000001000: n7538_o = n2110_o;
      13'b0000000000100: n7538_o = n5711_o;
      13'b0000000000010: n7538_o = n3260_o;
      13'b0000000000001: n7538_o = n2110_o;
      default: n7538_o = n2110_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7540_o = 1'b0;
      13'b0100000000000: n7540_o = n7350_o;
      13'b0010000000000: n7540_o = 1'b0;
      13'b0001000000000: n7540_o = 1'b0;
      13'b0000100000000: n7540_o = 1'b0;
      13'b0000010000000: n7540_o = 1'b0;
      13'b0000001000000: n7540_o = 1'b0;
      13'b0000000100000: n7540_o = 1'b0;
      13'b0000000010000: n7540_o = 1'b0;
      13'b0000000001000: n7540_o = n6016_o;
      13'b0000000000100: n7540_o = 1'b0;
      13'b0000000000010: n7540_o = 1'b0;
      13'b0000000000001: n7540_o = 1'b0;
      default: n7540_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7543_o = 1'b0;
      13'b0100000000000: n7543_o = n7352_o;
      13'b0010000000000: n7543_o = 1'b0;
      13'b0001000000000: n7543_o = 1'b0;
      13'b0000100000000: n7543_o = 1'b0;
      13'b0000010000000: n7543_o = 1'b0;
      13'b0000001000000: n7543_o = n6414_o;
      13'b0000000100000: n7543_o = 1'b0;
      13'b0000000010000: n7543_o = 1'b0;
      13'b0000000001000: n7543_o = n6017_o;
      13'b0000000000100: n7543_o = n5713_o;
      13'b0000000000010: n7543_o = 1'b0;
      13'b0000000000001: n7543_o = n3038_o;
      default: n7543_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7545_o = n1974_o;
      13'b0100000000000: n7545_o = n1974_o;
      13'b0010000000000: n7545_o = n1974_o;
      13'b0001000000000: n7545_o = n1974_o;
      13'b0000100000000: n7545_o = n1974_o;
      13'b0000010000000: n7545_o = n1974_o;
      13'b0000001000000: n7545_o = n1974_o;
      13'b0000000100000: n7545_o = n1974_o;
      13'b0000000010000: n7545_o = n6080_o;
      13'b0000000001000: n7545_o = n1974_o;
      13'b0000000000100: n7545_o = n5714_o;
      13'b0000000000010: n7545_o = n1974_o;
      13'b0000000000001: n7545_o = n1974_o;
      default: n7545_o = n1974_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7547_o = 1'b0;
      13'b0100000000000: n7547_o = 1'b0;
      13'b0010000000000: n7547_o = 1'b0;
      13'b0001000000000: n7547_o = 1'b0;
      13'b0000100000000: n7547_o = 1'b0;
      13'b0000010000000: n7547_o = 1'b0;
      13'b0000001000000: n7547_o = 1'b0;
      13'b0000000100000: n7547_o = 1'b0;
      13'b0000000010000: n7547_o = n6093_o;
      13'b0000000001000: n7547_o = 1'b0;
      13'b0000000000100: n7547_o = n5716_o;
      13'b0000000000010: n7547_o = 1'b0;
      13'b0000000000001: n7547_o = 1'b0;
      default: n7547_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7550_o = 1'b0;
      13'b0100000000000: n7550_o = 1'b0;
      13'b0010000000000: n7550_o = 1'b0;
      13'b0001000000000: n7550_o = 1'b0;
      13'b0000100000000: n7550_o = 1'b0;
      13'b0000010000000: n7550_o = 1'b0;
      13'b0000001000000: n7550_o = 1'b0;
      13'b0000000100000: n7550_o = 1'b0;
      13'b0000000010000: n7550_o = 1'b0;
      13'b0000000001000: n7550_o = 1'b0;
      13'b0000000000100: n7550_o = n5718_o;
      13'b0000000000010: n7550_o = 1'b0;
      13'b0000000000001: n7550_o = 1'b0;
      default: n7550_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7553_o = 1'b0;
      13'b0100000000000: n7553_o = n7354_o;
      13'b0010000000000: n7553_o = 1'b0;
      13'b0001000000000: n7553_o = 1'b0;
      13'b0000100000000: n7553_o = 1'b0;
      13'b0000010000000: n7553_o = 1'b0;
      13'b0000001000000: n7553_o = 1'b0;
      13'b0000000100000: n7553_o = 1'b0;
      13'b0000000010000: n7553_o = 1'b0;
      13'b0000000001000: n7553_o = 1'b0;
      13'b0000000000100: n7553_o = n5719_o;
      13'b0000000000010: n7553_o = 1'b0;
      13'b0000000000001: n7553_o = 1'b0;
      default: n7553_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7556_o = 1'b0;
      13'b0100000000000: n7556_o = 1'b0;
      13'b0010000000000: n7556_o = n7007_o;
      13'b0001000000000: n7556_o = n6748_o;
      13'b0000100000000: n7556_o = 1'b0;
      13'b0000010000000: n7556_o = n6532_o;
      13'b0000001000000: n7556_o = 1'b0;
      13'b0000000100000: n7556_o = 1'b0;
      13'b0000000010000: n7556_o = 1'b0;
      13'b0000000001000: n7556_o = 1'b0;
      13'b0000000000100: n7556_o = n5720_o;
      13'b0000000000010: n7556_o = n3273_o;
      13'b0000000000001: n7556_o = 1'b0;
      default: n7556_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7559_o = 1'b0;
      13'b0100000000000: n7559_o = n7356_o;
      13'b0010000000000: n7559_o = n7009_o;
      13'b0001000000000: n7559_o = n6750_o;
      13'b0000100000000: n7559_o = 1'b0;
      13'b0000010000000: n7559_o = n6534_o;
      13'b0000001000000: n7559_o = n6415_o;
      13'b0000000100000: n7559_o = 1'b0;
      13'b0000000010000: n7559_o = 1'b0;
      13'b0000000001000: n7559_o = 1'b0;
      13'b0000000000100: n7559_o = n5721_o;
      13'b0000000000010: n7559_o = n3276_o;
      13'b0000000000001: n7559_o = 1'b0;
      default: n7559_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7562_o = 1'b0;
      13'b0100000000000: n7562_o = n7358_o;
      13'b0010000000000: n7562_o = 1'b0;
      13'b0001000000000: n7562_o = 1'b0;
      13'b0000100000000: n7562_o = 1'b0;
      13'b0000010000000: n7562_o = 1'b0;
      13'b0000001000000: n7562_o = 1'b0;
      13'b0000000100000: n7562_o = 1'b0;
      13'b0000000010000: n7562_o = 1'b0;
      13'b0000000001000: n7562_o = 1'b0;
      13'b0000000000100: n7562_o = 1'b0;
      13'b0000000000010: n7562_o = 1'b0;
      13'b0000000000001: n7562_o = 1'b0;
      default: n7562_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7565_o = 1'b0;
      13'b0100000000000: n7565_o = n7360_o;
      13'b0010000000000: n7565_o = 1'b0;
      13'b0001000000000: n7565_o = 1'b0;
      13'b0000100000000: n7565_o = 1'b0;
      13'b0000010000000: n7565_o = 1'b0;
      13'b0000001000000: n7565_o = 1'b0;
      13'b0000000100000: n7565_o = 1'b0;
      13'b0000000010000: n7565_o = 1'b0;
      13'b0000000001000: n7565_o = 1'b0;
      13'b0000000000100: n7565_o = n5723_o;
      13'b0000000000010: n7565_o = 1'b0;
      13'b0000000000001: n7565_o = n3040_o;
      default: n7565_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7568_o = 1'b0;
      13'b0100000000000: n7568_o = 1'b0;
      13'b0010000000000: n7568_o = n7011_o;
      13'b0001000000000: n7568_o = n6752_o;
      13'b0000100000000: n7568_o = 1'b0;
      13'b0000010000000: n7568_o = n6536_o;
      13'b0000001000000: n7568_o = 1'b0;
      13'b0000000100000: n7568_o = 1'b0;
      13'b0000000010000: n7568_o = 1'b0;
      13'b0000000001000: n7568_o = 1'b0;
      13'b0000000000100: n7568_o = n5725_o;
      13'b0000000000010: n7568_o = n3278_o;
      13'b0000000000001: n7568_o = 1'b0;
      default: n7568_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7571_o = 1'b0;
      13'b0100000000000: n7571_o = n7362_o;
      13'b0010000000000: n7571_o = 1'b0;
      13'b0001000000000: n7571_o = 1'b0;
      13'b0000100000000: n7571_o = 1'b0;
      13'b0000010000000: n7571_o = 1'b0;
      13'b0000001000000: n7571_o = 1'b0;
      13'b0000000100000: n7571_o = 1'b0;
      13'b0000000010000: n7571_o = 1'b0;
      13'b0000000001000: n7571_o = 1'b0;
      13'b0000000000100: n7571_o = n5727_o;
      13'b0000000000010: n7571_o = 1'b0;
      13'b0000000000001: n7571_o = 1'b0;
      default: n7571_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7574_o = 1'b0;
      13'b0100000000000: n7574_o = 1'b0;
      13'b0010000000000: n7574_o = n7012_o;
      13'b0001000000000: n7574_o = n6754_o;
      13'b0000100000000: n7574_o = 1'b0;
      13'b0000010000000: n7574_o = n6538_o;
      13'b0000001000000: n7574_o = n6416_o;
      13'b0000000100000: n7574_o = n6111_o;
      13'b0000000010000: n7574_o = 1'b0;
      13'b0000000001000: n7574_o = 1'b0;
      13'b0000000000100: n7574_o = n5728_o;
      13'b0000000000010: n7574_o = n3280_o;
      13'b0000000000001: n7574_o = n3042_o;
      default: n7574_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7576_o = n1861_o;
      13'b0100000000000: n7576_o = n7065_o;
      13'b0010000000000: n7576_o = n1861_o;
      13'b0001000000000: n7576_o = n1861_o;
      13'b0000100000000: n7576_o = n1861_o;
      13'b0000010000000: n7576_o = n1861_o;
      13'b0000001000000: n7576_o = n1861_o;
      13'b0000000100000: n7576_o = n1861_o;
      13'b0000000010000: n7576_o = n1861_o;
      13'b0000000001000: n7576_o = n1861_o;
      13'b0000000000100: n7576_o = n1861_o;
      13'b0000000000010: n7576_o = n1861_o;
      13'b0000000000001: n7576_o = n1861_o;
      default: n7576_o = n1861_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7577_o = n1867_o;
      13'b0100000000000: n7577_o = n1867_o;
      13'b0010000000000: n7577_o = n1867_o;
      13'b0001000000000: n7577_o = n1867_o;
      13'b0000100000000: n7577_o = n1867_o;
      13'b0000010000000: n7577_o = n1867_o;
      13'b0000001000000: n7577_o = n1867_o;
      13'b0000000100000: n7577_o = n1867_o;
      13'b0000000010000: n7577_o = n1867_o;
      13'b0000000001000: n7577_o = n1867_o;
      13'b0000000000100: n7577_o = n5729_o;
      13'b0000000000010: n7577_o = n1867_o;
      13'b0000000000001: n7577_o = n1867_o;
      default: n7577_o = n1867_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7579_o = 1'b0;
      13'b0100000000000: n7579_o = 1'b0;
      13'b0010000000000: n7579_o = 1'b0;
      13'b0001000000000: n7579_o = 1'b0;
      13'b0000100000000: n7579_o = 1'b0;
      13'b0000010000000: n7579_o = 1'b0;
      13'b0000001000000: n7579_o = 1'b0;
      13'b0000000100000: n7579_o = 1'b0;
      13'b0000000010000: n7579_o = 1'b0;
      13'b0000000001000: n7579_o = 1'b0;
      13'b0000000000100: n7579_o = n5731_o;
      13'b0000000000010: n7579_o = 1'b0;
      13'b0000000000001: n7579_o = 1'b0;
      default: n7579_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7581_o = n2113_o;
      13'b0100000000000: n7581_o = n2113_o;
      13'b0010000000000: n7581_o = n2113_o;
      13'b0001000000000: n7581_o = n2113_o;
      13'b0000100000000: n7581_o = n2113_o;
      13'b0000010000000: n7581_o = n2113_o;
      13'b0000001000000: n7581_o = n6417_o;
      13'b0000000100000: n7581_o = n2113_o;
      13'b0000000010000: n7581_o = n2113_o;
      13'b0000000001000: n7581_o = n2113_o;
      13'b0000000000100: n7581_o = n5732_o;
      13'b0000000000010: n7581_o = n2113_o;
      13'b0000000000001: n7581_o = n3043_o;
      default: n7581_o = n2113_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7584_o = n7523_o;
      13'b0100000000000: n7584_o = n7365_o;
      13'b0010000000000: n7584_o = n7013_o;
      13'b0001000000000: n7584_o = n6755_o;
      13'b0000100000000: n7584_o = 1'b0;
      13'b0000010000000: n7584_o = n6541_o;
      13'b0000001000000: n7584_o = n6418_o;
      13'b0000000100000: n7584_o = n6114_o;
      13'b0000000010000: n7584_o = 1'b0;
      13'b0000000001000: n7584_o = n6018_o;
      13'b0000000000100: n7584_o = n5733_o;
      13'b0000000000010: n7584_o = n3283_o;
      13'b0000000000001: n7584_o = n3045_o;
      default: n7584_o = 1'b1;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7587_o = n7524_o;
      13'b0100000000000: n7587_o = 1'b0;
      13'b0010000000000: n7587_o = 1'b0;
      13'b0001000000000: n7587_o = 1'b0;
      13'b0000100000000: n7587_o = 1'b0;
      13'b0000010000000: n7587_o = 1'b0;
      13'b0000001000000: n7587_o = 1'b0;
      13'b0000000100000: n7587_o = 1'b0;
      13'b0000000010000: n7587_o = 1'b0;
      13'b0000000001000: n7587_o = 1'b0;
      13'b0000000000100: n7587_o = n5735_o;
      13'b0000000000010: n7587_o = 1'b0;
      13'b0000000000001: n7587_o = n3047_o;
      default: n7587_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7591_o = 1'b0;
      13'b0100000000000: n7591_o = 1'b0;
      13'b0010000000000: n7591_o = 1'b0;
      13'b0001000000000: n7591_o = 1'b0;
      13'b0000100000000: n7591_o = 1'b1;
      13'b0000010000000: n7591_o = 1'b0;
      13'b0000001000000: n7591_o = 1'b0;
      13'b0000000100000: n7591_o = 1'b0;
      13'b0000000010000: n7591_o = 1'b0;
      13'b0000000001000: n7591_o = 1'b0;
      13'b0000000000100: n7591_o = 1'b0;
      13'b0000000000010: n7591_o = 1'b0;
      13'b0000000000001: n7591_o = 1'b0;
      default: n7591_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7594_o = n7525_o;
      13'b0100000000000: n7594_o = 1'b0;
      13'b0010000000000: n7594_o = 1'b0;
      13'b0001000000000: n7594_o = 1'b0;
      13'b0000100000000: n7594_o = 1'b0;
      13'b0000010000000: n7594_o = 1'b0;
      13'b0000001000000: n7594_o = 1'b0;
      13'b0000000100000: n7594_o = 1'b0;
      13'b0000000010000: n7594_o = 1'b0;
      13'b0000000001000: n7594_o = 1'b0;
      13'b0000000000100: n7594_o = 1'b0;
      13'b0000000000010: n7594_o = 1'b0;
      13'b0000000000001: n7594_o = 1'b0;
      default: n7594_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7597_o = 1'b0;
      13'b0100000000000: n7597_o = 1'b0;
      13'b0010000000000: n7597_o = 1'b0;
      13'b0001000000000: n7597_o = 1'b0;
      13'b0000100000000: n7597_o = 1'b0;
      13'b0000010000000: n7597_o = 1'b0;
      13'b0000001000000: n7597_o = 1'b0;
      13'b0000000100000: n7597_o = 1'b0;
      13'b0000000010000: n7597_o = 1'b0;
      13'b0000000001000: n7597_o = 1'b0;
      13'b0000000000100: n7597_o = n5737_o;
      13'b0000000000010: n7597_o = 1'b0;
      13'b0000000000001: n7597_o = 1'b0;
      default: n7597_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7600_o = 1'b0;
      13'b0100000000000: n7600_o = 1'b0;
      13'b0010000000000: n7600_o = 1'b0;
      13'b0001000000000: n7600_o = 1'b0;
      13'b0000100000000: n7600_o = 1'b0;
      13'b0000010000000: n7600_o = 1'b0;
      13'b0000001000000: n7600_o = 1'b0;
      13'b0000000100000: n7600_o = 1'b0;
      13'b0000000010000: n7600_o = 1'b0;
      13'b0000000001000: n7600_o = n6020_o;
      13'b0000000000100: n7600_o = n5739_o;
      13'b0000000000010: n7600_o = 1'b0;
      13'b0000000000001: n7600_o = 1'b0;
      default: n7600_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7606_o = 1'b1;
      13'b0100000000000: n7606_o = n7367_o;
      13'b0010000000000: n7606_o = n7014_o;
      13'b0001000000000: n7606_o = n6756_o;
      13'b0000100000000: n7606_o = 1'b1;
      13'b0000010000000: n7606_o = n6544_o;
      13'b0000001000000: n7606_o = n6419_o;
      13'b0000000100000: n7606_o = n6117_o;
      13'b0000000010000: n7606_o = 1'b0;
      13'b0000000001000: n7606_o = n6021_o;
      13'b0000000000100: n7606_o = n5740_o;
      13'b0000000000010: n7606_o = n3286_o;
      13'b0000000000001: n7606_o = n3049_o;
      default: n7606_o = 1'b1;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7609_o = 1'b0;
      13'b0100000000000: n7609_o = 1'b0;
      13'b0010000000000: n7609_o = 1'b0;
      13'b0001000000000: n7609_o = 1'b0;
      13'b0000100000000: n7609_o = 1'b0;
      13'b0000010000000: n7609_o = 1'b0;
      13'b0000001000000: n7609_o = 1'b0;
      13'b0000000100000: n7609_o = 1'b0;
      13'b0000000010000: n7609_o = 1'b0;
      13'b0000000001000: n7609_o = 1'b0;
      13'b0000000000100: n7609_o = n5742_o;
      13'b0000000000010: n7609_o = 1'b0;
      13'b0000000000001: n7609_o = 1'b0;
      default: n7609_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7612_o = 1'b0;
      13'b0100000000000: n7612_o = n7369_o;
      13'b0010000000000: n7612_o = n7016_o;
      13'b0001000000000: n7612_o = n6757_o;
      13'b0000100000000: n7612_o = 1'b0;
      13'b0000010000000: n7612_o = n6547_o;
      13'b0000001000000: n7612_o = n6421_o;
      13'b0000000100000: n7612_o = 1'b0;
      13'b0000000010000: n7612_o = 1'b0;
      13'b0000000001000: n7612_o = n6022_o;
      13'b0000000000100: n7612_o = n5743_o;
      13'b0000000000010: n7612_o = n3289_o;
      13'b0000000000001: n7612_o = n3051_o;
      default: n7612_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7615_o = 1'b0;
      13'b0100000000000: n7615_o = 1'b0;
      13'b0010000000000: n7615_o = n7018_o;
      13'b0001000000000: n7615_o = n6759_o;
      13'b0000100000000: n7615_o = 1'b0;
      13'b0000010000000: n7615_o = n6549_o;
      13'b0000001000000: n7615_o = n6423_o;
      13'b0000000100000: n7615_o = 1'b0;
      13'b0000000010000: n7615_o = 1'b0;
      13'b0000000001000: n7615_o = 1'b0;
      13'b0000000000100: n7615_o = 1'b0;
      13'b0000000000010: n7615_o = 1'b0;
      13'b0000000000001: n7615_o = 1'b0;
      default: n7615_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7618_o = 1'b0;
      13'b0100000000000: n7618_o = 1'b0;
      13'b0010000000000: n7618_o = n7020_o;
      13'b0001000000000: n7618_o = 1'b0;
      13'b0000100000000: n7618_o = 1'b0;
      13'b0000010000000: n7618_o = n6551_o;
      13'b0000001000000: n7618_o = n6425_o;
      13'b0000000100000: n7618_o = 1'b0;
      13'b0000000010000: n7618_o = 1'b0;
      13'b0000000001000: n7618_o = 1'b0;
      13'b0000000000100: n7618_o = 1'b0;
      13'b0000000000010: n7618_o = 1'b0;
      13'b0000000000001: n7618_o = 1'b0;
      default: n7618_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7621_o = 1'b0;
      13'b0100000000000: n7621_o = 1'b0;
      13'b0010000000000: n7621_o = 1'b0;
      13'b0001000000000: n7621_o = 1'b0;
      13'b0000100000000: n7621_o = 1'b0;
      13'b0000010000000: n7621_o = 1'b0;
      13'b0000001000000: n7621_o = 1'b0;
      13'b0000000100000: n7621_o = 1'b0;
      13'b0000000010000: n7621_o = 1'b0;
      13'b0000000001000: n7621_o = 1'b0;
      13'b0000000000100: n7621_o = 1'b0;
      13'b0000000000010: n7621_o = 1'b0;
      13'b0000000000001: n7621_o = n3053_o;
      default: n7621_o = 1'b0;
    endcase
  assign n7623_o = n1870_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7624_o = n7623_o;
      13'b0100000000000: n7624_o = n7623_o;
      13'b0010000000000: n7624_o = n7623_o;
      13'b0001000000000: n7624_o = n7623_o;
      13'b0000100000000: n7624_o = n7623_o;
      13'b0000010000000: n7624_o = n7623_o;
      13'b0000001000000: n7624_o = n7623_o;
      13'b0000000100000: n7624_o = n7623_o;
      13'b0000000010000: n7624_o = n7623_o;
      13'b0000000001000: n7624_o = n7623_o;
      13'b0000000000100: n7624_o = n5749_o;
      13'b0000000000010: n7624_o = n7623_o;
      13'b0000000000001: n7624_o = n7623_o;
      default: n7624_o = n7623_o;
    endcase
  assign n7625_o = n1870_o[19:17];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7626_o = n7625_o;
      13'b0100000000000: n7626_o = n7625_o;
      13'b0010000000000: n7626_o = n7625_o;
      13'b0001000000000: n7626_o = n7625_o;
      13'b0000100000000: n7626_o = n7625_o;
      13'b0000010000000: n7626_o = n7625_o;
      13'b0000001000000: n7626_o = n7625_o;
      13'b0000000100000: n7626_o = n7625_o;
      13'b0000000010000: n7626_o = n7625_o;
      13'b0000000001000: n7626_o = n7625_o;
      13'b0000000000100: n7626_o = n7625_o;
      13'b0000000000010: n7626_o = n7625_o;
      13'b0000000000001: n7626_o = n3057_o;
      default: n7626_o = n7625_o;
    endcase
  assign n7627_o = n1870_o[20];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7628_o = n7627_o;
      13'b0100000000000: n7628_o = n7627_o;
      13'b0010000000000: n7628_o = n7627_o;
      13'b0001000000000: n7628_o = n7627_o;
      13'b0000100000000: n7628_o = n7627_o;
      13'b0000010000000: n7628_o = n7627_o;
      13'b0000001000000: n7628_o = n7627_o;
      13'b0000000100000: n7628_o = n7627_o;
      13'b0000000010000: n7628_o = n7627_o;
      13'b0000000001000: n7628_o = n7627_o;
      13'b0000000000100: n7628_o = n5751_o;
      13'b0000000000010: n7628_o = n7627_o;
      13'b0000000000001: n7628_o = n7627_o;
      default: n7628_o = n7627_o;
    endcase
  assign n7629_o = n1870_o[24];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7630_o = n7629_o;
      13'b0100000000000: n7630_o = n7629_o;
      13'b0010000000000: n7630_o = n7629_o;
      13'b0001000000000: n7630_o = n7629_o;
      13'b0000100000000: n7630_o = n7629_o;
      13'b0000010000000: n7630_o = n7629_o;
      13'b0000001000000: n7630_o = n7629_o;
      13'b0000000100000: n7630_o = n7629_o;
      13'b0000000010000: n7630_o = n7629_o;
      13'b0000000001000: n7630_o = n7629_o;
      13'b0000000000100: n7630_o = n5753_o;
      13'b0000000000010: n7630_o = n7629_o;
      13'b0000000000001: n7630_o = n7629_o;
      default: n7630_o = n7629_o;
    endcase
  assign n7631_o = n1870_o[26];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7632_o = n7631_o;
      13'b0100000000000: n7632_o = n7631_o;
      13'b0010000000000: n7632_o = n7631_o;
      13'b0001000000000: n7632_o = n7631_o;
      13'b0000100000000: n7632_o = n7631_o;
      13'b0000010000000: n7632_o = n7631_o;
      13'b0000001000000: n7632_o = n7631_o;
      13'b0000000100000: n7632_o = n7631_o;
      13'b0000000010000: n7632_o = n7631_o;
      13'b0000000001000: n7632_o = n7631_o;
      13'b0000000000100: n7632_o = n7631_o;
      13'b0000000000010: n7632_o = n7631_o;
      13'b0000000000001: n7632_o = n3059_o;
      default: n7632_o = n7631_o;
    endcase
  assign n7633_o = n1870_o[29];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7634_o = n7633_o;
      13'b0100000000000: n7634_o = n7371_o;
      13'b0010000000000: n7634_o = n7633_o;
      13'b0001000000000: n7634_o = n7633_o;
      13'b0000100000000: n7634_o = n7633_o;
      13'b0000010000000: n7634_o = n7633_o;
      13'b0000001000000: n7634_o = n7633_o;
      13'b0000000100000: n7634_o = n7633_o;
      13'b0000000010000: n7634_o = n7633_o;
      13'b0000000001000: n7634_o = n7633_o;
      13'b0000000000100: n7634_o = n7633_o;
      13'b0000000000010: n7634_o = n7633_o;
      13'b0000000000001: n7634_o = n7633_o;
      default: n7634_o = n7633_o;
    endcase
  assign n7635_o = n1870_o[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7636_o = n7635_o;
      13'b0100000000000: n7636_o = n7635_o;
      13'b0010000000000: n7636_o = n7022_o;
      13'b0001000000000: n7636_o = n7635_o;
      13'b0000100000000: n7636_o = n7635_o;
      13'b0000010000000: n7636_o = n7635_o;
      13'b0000001000000: n7636_o = n7635_o;
      13'b0000000100000: n7636_o = n7635_o;
      13'b0000000010000: n7636_o = n7635_o;
      13'b0000000001000: n7636_o = n7635_o;
      13'b0000000000100: n7636_o = n5755_o;
      13'b0000000000010: n7636_o = n7635_o;
      13'b0000000000001: n7636_o = n7635_o;
      default: n7636_o = n7635_o;
    endcase
  assign n7637_o = n1870_o[36];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7638_o = n7637_o;
      13'b0100000000000: n7638_o = n7637_o;
      13'b0010000000000: n7638_o = n7637_o;
      13'b0001000000000: n7638_o = n7637_o;
      13'b0000100000000: n7638_o = n7637_o;
      13'b0000010000000: n7638_o = n7637_o;
      13'b0000001000000: n7638_o = n7637_o;
      13'b0000000100000: n7638_o = n7637_o;
      13'b0000000010000: n7638_o = n7637_o;
      13'b0000000001000: n7638_o = n7637_o;
      13'b0000000000100: n7638_o = n5757_o;
      13'b0000000000010: n7638_o = n7637_o;
      13'b0000000000001: n7638_o = n7637_o;
      default: n7638_o = n7637_o;
    endcase
  assign n7639_o = n1870_o[37];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7640_o = n7639_o;
      13'b0100000000000: n7640_o = n7639_o;
      13'b0010000000000: n7640_o = n7639_o;
      13'b0001000000000: n7640_o = n7639_o;
      13'b0000100000000: n7640_o = n7639_o;
      13'b0000010000000: n7640_o = n7639_o;
      13'b0000001000000: n7640_o = n7639_o;
      13'b0000000100000: n7640_o = n7639_o;
      13'b0000000010000: n7640_o = n7639_o;
      13'b0000000001000: n7640_o = n7639_o;
      13'b0000000000100: n7640_o = n7639_o;
      13'b0000000000010: n7640_o = n7639_o;
      13'b0000000000001: n7640_o = n3061_o;
      default: n7640_o = n7639_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7641_o = n1966_o;
      13'b0100000000000: n7641_o = n1966_o;
      13'b0010000000000: n7641_o = n1966_o;
      13'b0001000000000: n7641_o = n6760_o;
      13'b0000100000000: n7641_o = n1966_o;
      13'b0000010000000: n7641_o = n1966_o;
      13'b0000001000000: n7641_o = n1966_o;
      13'b0000000100000: n7641_o = n1966_o;
      13'b0000000010000: n7641_o = n1966_o;
      13'b0000000001000: n7641_o = n1966_o;
      13'b0000000000100: n7641_o = n1966_o;
      13'b0000000000010: n7641_o = n1966_o;
      13'b0000000000001: n7641_o = n1966_o;
      default: n7641_o = n1966_o;
    endcase
  assign n7642_o = n1870_o[39];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7643_o = n7642_o;
      13'b0100000000000: n7643_o = n7642_o;
      13'b0010000000000: n7643_o = n7642_o;
      13'b0001000000000: n7643_o = n7642_o;
      13'b0000100000000: n7643_o = n7642_o;
      13'b0000010000000: n7643_o = n7642_o;
      13'b0000001000000: n7643_o = n7642_o;
      13'b0000000100000: n7643_o = n7642_o;
      13'b0000000010000: n7643_o = n7642_o;
      13'b0000000001000: n7643_o = n7642_o;
      13'b0000000000100: n7643_o = n7642_o;
      13'b0000000000010: n7643_o = n7642_o;
      13'b0000000000001: n7643_o = n3063_o;
      default: n7643_o = n7642_o;
    endcase
  assign n7644_o = n1870_o[40];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7645_o = n7644_o;
      13'b0100000000000: n7645_o = n7644_o;
      13'b0010000000000: n7645_o = n7644_o;
      13'b0001000000000: n7645_o = n7644_o;
      13'b0000100000000: n7645_o = n7644_o;
      13'b0000010000000: n7645_o = n7644_o;
      13'b0000001000000: n7645_o = n7644_o;
      13'b0000000100000: n7645_o = n7644_o;
      13'b0000000010000: n7645_o = n7644_o;
      13'b0000000001000: n7645_o = n7644_o;
      13'b0000000000100: n7645_o = n5759_o;
      13'b0000000000010: n7645_o = n3263_o;
      13'b0000000000001: n7645_o = n7644_o;
      default: n7645_o = n7644_o;
    endcase
  assign n7646_o = n3065_o[0];
  assign n7647_o = n1870_o[42];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7648_o = n7647_o;
      13'b0100000000000: n7648_o = n7373_o;
      13'b0010000000000: n7648_o = n7647_o;
      13'b0001000000000: n7648_o = n7647_o;
      13'b0000100000000: n7648_o = n7647_o;
      13'b0000010000000: n7648_o = n7647_o;
      13'b0000001000000: n7648_o = n7647_o;
      13'b0000000100000: n7648_o = n7647_o;
      13'b0000000010000: n7648_o = n7647_o;
      13'b0000000001000: n7648_o = n7647_o;
      13'b0000000000100: n7648_o = n5761_o;
      13'b0000000000010: n7648_o = n7647_o;
      13'b0000000000001: n7648_o = n7646_o;
      default: n7648_o = n7647_o;
    endcase
  assign n7649_o = n3065_o[1];
  assign n7650_o = n1870_o[43];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7651_o = n7650_o;
      13'b0100000000000: n7651_o = n7650_o;
      13'b0010000000000: n7651_o = n7650_o;
      13'b0001000000000: n7651_o = n7650_o;
      13'b0000100000000: n7651_o = n7650_o;
      13'b0000010000000: n7651_o = n7650_o;
      13'b0000001000000: n7651_o = n7650_o;
      13'b0000000100000: n7651_o = n7650_o;
      13'b0000000010000: n7651_o = n7650_o;
      13'b0000000001000: n7651_o = n7650_o;
      13'b0000000000100: n7651_o = n5763_o;
      13'b0000000000010: n7651_o = n7650_o;
      13'b0000000000001: n7651_o = n7649_o;
      default: n7651_o = n7650_o;
    endcase
  assign n7652_o = n1870_o[44];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7653_o = n7652_o;
      13'b0100000000000: n7653_o = n7652_o;
      13'b0010000000000: n7653_o = n7652_o;
      13'b0001000000000: n7653_o = n7652_o;
      13'b0000100000000: n7653_o = n7652_o;
      13'b0000010000000: n7653_o = n7652_o;
      13'b0000001000000: n7653_o = n6427_o;
      13'b0000000100000: n7653_o = n7652_o;
      13'b0000000010000: n7653_o = n7652_o;
      13'b0000000001000: n7653_o = n7652_o;
      13'b0000000000100: n7653_o = n5765_o;
      13'b0000000000010: n7653_o = n7652_o;
      13'b0000000000001: n7653_o = n7652_o;
      default: n7653_o = n7652_o;
    endcase
  assign n7654_o = n3264_o[0];
  assign n7655_o = n5769_o[0];
  assign n7656_o = n2121_o[0];
  assign n7657_o = n1870_o[46];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n7658_o = n1996_o ? n7656_o : n7657_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7659_o = n7658_o;
      13'b0100000000000: n7659_o = n7658_o;
      13'b0010000000000: n7659_o = n7658_o;
      13'b0001000000000: n7659_o = n6764_o;
      13'b0000100000000: n7659_o = n7658_o;
      13'b0000010000000: n7659_o = n7658_o;
      13'b0000001000000: n7659_o = n7658_o;
      13'b0000000100000: n7659_o = n7658_o;
      13'b0000000010000: n7659_o = n7658_o;
      13'b0000000001000: n7659_o = n7658_o;
      13'b0000000000100: n7659_o = n7655_o;
      13'b0000000000010: n7659_o = n7654_o;
      13'b0000000000001: n7659_o = n7658_o;
      default: n7659_o = n7658_o;
    endcase
  assign n7660_o = n3264_o[1];
  assign n7661_o = n5769_o[1];
  assign n7662_o = n2121_o[1];
  assign n7663_o = n1870_o[47];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1586:17  */
  assign n7664_o = n1996_o ? n7662_o : n7663_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7665_o = n7664_o;
      13'b0100000000000: n7665_o = n7664_o;
      13'b0010000000000: n7665_o = n7664_o;
      13'b0001000000000: n7665_o = n7664_o;
      13'b0000100000000: n7665_o = n7664_o;
      13'b0000010000000: n7665_o = n7664_o;
      13'b0000001000000: n7665_o = n7664_o;
      13'b0000000100000: n7665_o = n7664_o;
      13'b0000000010000: n7665_o = n6097_o;
      13'b0000000001000: n7665_o = n7664_o;
      13'b0000000000100: n7665_o = n7661_o;
      13'b0000000000010: n7665_o = n7660_o;
      13'b0000000000001: n7665_o = n7664_o;
      default: n7665_o = n7664_o;
    endcase
  assign n7666_o = n5769_o[2];
  assign n7667_o = n1870_o[48];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7668_o = n7667_o;
      13'b0100000000000: n7668_o = n7667_o;
      13'b0010000000000: n7668_o = n7667_o;
      13'b0001000000000: n7668_o = n7667_o;
      13'b0000100000000: n7668_o = n7667_o;
      13'b0000010000000: n7668_o = n7667_o;
      13'b0000001000000: n7668_o = n7667_o;
      13'b0000000100000: n7668_o = n7667_o;
      13'b0000000010000: n7668_o = n7667_o;
      13'b0000000001000: n7668_o = n7667_o;
      13'b0000000000100: n7668_o = n7666_o;
      13'b0000000000010: n7668_o = n7667_o;
      13'b0000000000001: n7668_o = n7667_o;
      default: n7668_o = n7667_o;
    endcase
  assign n7669_o = n3296_o[0];
  assign n7670_o = n1870_o[49];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7671_o = n7670_o;
      13'b0100000000000: n7671_o = n7670_o;
      13'b0010000000000: n7671_o = n7670_o;
      13'b0001000000000: n7671_o = n7670_o;
      13'b0000100000000: n7671_o = n7670_o;
      13'b0000010000000: n7671_o = n6527_o;
      13'b0000001000000: n7671_o = n6429_o;
      13'b0000000100000: n7671_o = n7670_o;
      13'b0000000010000: n7671_o = n7670_o;
      13'b0000000001000: n7671_o = n6024_o;
      13'b0000000000100: n7671_o = n5771_o;
      13'b0000000000010: n7671_o = n7669_o;
      13'b0000000000001: n7671_o = n3067_o;
      default: n7671_o = n7670_o;
    endcase
  assign n7672_o = n3296_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7673_o = n2127_o;
      13'b0100000000000: n7673_o = n2127_o;
      13'b0010000000000: n7673_o = n2127_o;
      13'b0001000000000: n7673_o = n6765_o;
      13'b0000100000000: n7673_o = n2127_o;
      13'b0000010000000: n7673_o = n2127_o;
      13'b0000001000000: n7673_o = n2127_o;
      13'b0000000100000: n7673_o = n2127_o;
      13'b0000000010000: n7673_o = n2127_o;
      13'b0000000001000: n7673_o = n2127_o;
      13'b0000000000100: n7673_o = n2127_o;
      13'b0000000000010: n7673_o = n7672_o;
      13'b0000000000001: n7673_o = n3069_o;
      default: n7673_o = n2127_o;
    endcase
  assign n7674_o = n5774_o[1:0];
  assign n7675_o = n1870_o[52:51];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7676_o = n7675_o;
      13'b0100000000000: n7676_o = n7675_o;
      13'b0010000000000: n7676_o = n7675_o;
      13'b0001000000000: n7676_o = n7675_o;
      13'b0000100000000: n7676_o = n7675_o;
      13'b0000010000000: n7676_o = n7675_o;
      13'b0000001000000: n7676_o = n7675_o;
      13'b0000000100000: n7676_o = n7675_o;
      13'b0000000010000: n7676_o = n7675_o;
      13'b0000000001000: n7676_o = n7675_o;
      13'b0000000000100: n7676_o = n7674_o;
      13'b0000000000010: n7676_o = n7675_o;
      13'b0000000000001: n7676_o = n3071_o;
      default: n7676_o = n7675_o;
    endcase
  assign n7677_o = n5774_o[2];
  assign n7678_o = n1870_o[53];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7679_o = n7678_o;
      13'b0100000000000: n7679_o = n7678_o;
      13'b0010000000000: n7679_o = n7678_o;
      13'b0001000000000: n7679_o = n7678_o;
      13'b0000100000000: n7679_o = n7678_o;
      13'b0000010000000: n7679_o = n7678_o;
      13'b0000001000000: n7679_o = n7678_o;
      13'b0000000100000: n7679_o = n7678_o;
      13'b0000000010000: n7679_o = n7678_o;
      13'b0000000001000: n7679_o = n5831_o;
      13'b0000000000100: n7679_o = n7677_o;
      13'b0000000000010: n7679_o = n7678_o;
      13'b0000000000001: n7679_o = n7678_o;
      default: n7679_o = n7678_o;
    endcase
  assign n7680_o = n5774_o[3];
  assign n7681_o = n1870_o[54];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7682_o = n7681_o;
      13'b0100000000000: n7682_o = n7681_o;
      13'b0010000000000: n7682_o = n7681_o;
      13'b0001000000000: n7682_o = n7681_o;
      13'b0000100000000: n7682_o = n7681_o;
      13'b0000010000000: n7682_o = n7681_o;
      13'b0000001000000: n7682_o = n7681_o;
      13'b0000000100000: n7682_o = n7681_o;
      13'b0000000010000: n7682_o = n7681_o;
      13'b0000000001000: n7682_o = n7681_o;
      13'b0000000000100: n7682_o = n7680_o;
      13'b0000000000010: n7682_o = n7681_o;
      13'b0000000000001: n7682_o = n7681_o;
      default: n7682_o = n7681_o;
    endcase
  assign n7683_o = n3073_o[0];
  assign n7684_o = n5774_o[4];
  assign n7685_o = n1870_o[55];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7686_o = n7685_o;
      13'b0100000000000: n7686_o = n7375_o;
      13'b0010000000000: n7686_o = n7685_o;
      13'b0001000000000: n7686_o = n7685_o;
      13'b0000100000000: n7686_o = n7685_o;
      13'b0000010000000: n7686_o = n7685_o;
      13'b0000001000000: n7686_o = n7685_o;
      13'b0000000100000: n7686_o = n7685_o;
      13'b0000000010000: n7686_o = n7685_o;
      13'b0000000001000: n7686_o = n7685_o;
      13'b0000000000100: n7686_o = n7684_o;
      13'b0000000000010: n7686_o = n7685_o;
      13'b0000000000001: n7686_o = n7683_o;
      default: n7686_o = n7685_o;
    endcase
  assign n7687_o = n3073_o[1];
  assign n7688_o = n1870_o[56];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7689_o = n7688_o;
      13'b0100000000000: n7689_o = n7688_o;
      13'b0010000000000: n7689_o = n7688_o;
      13'b0001000000000: n7689_o = n6766_o;
      13'b0000100000000: n7689_o = n7688_o;
      13'b0000010000000: n7689_o = n6481_o;
      13'b0000001000000: n7689_o = n6431_o;
      13'b0000000100000: n7689_o = n7688_o;
      13'b0000000010000: n7689_o = n7688_o;
      13'b0000000001000: n7689_o = n6028_o;
      13'b0000000000100: n7689_o = n5776_o;
      13'b0000000000010: n7689_o = n7688_o;
      13'b0000000000001: n7689_o = n7687_o;
      default: n7689_o = n7688_o;
    endcase
  assign n7690_o = n1870_o[60:57];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7691_o = n7690_o;
      13'b0100000000000: n7691_o = n7690_o;
      13'b0010000000000: n7691_o = n7690_o;
      13'b0001000000000: n7691_o = n7690_o;
      13'b0000100000000: n7691_o = n7690_o;
      13'b0000010000000: n7691_o = n7690_o;
      13'b0000001000000: n7691_o = n7690_o;
      13'b0000000100000: n7691_o = n7690_o;
      13'b0000000010000: n7691_o = n7690_o;
      13'b0000000001000: n7691_o = n7690_o;
      13'b0000000000100: n7691_o = n5779_o;
      13'b0000000000010: n7691_o = n7690_o;
      13'b0000000000001: n7691_o = n7690_o;
      default: n7691_o = n7690_o;
    endcase
  assign n7692_o = n1870_o[61];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7693_o = n7692_o;
      13'b0100000000000: n7693_o = n7692_o;
      13'b0010000000000: n7693_o = n7024_o;
      13'b0001000000000: n7693_o = n7692_o;
      13'b0000100000000: n7693_o = n7692_o;
      13'b0000010000000: n7693_o = n7692_o;
      13'b0000001000000: n7693_o = n7692_o;
      13'b0000000100000: n7693_o = n7692_o;
      13'b0000000010000: n7693_o = n7692_o;
      13'b0000000001000: n7693_o = n7692_o;
      13'b0000000000100: n7693_o = n7692_o;
      13'b0000000000010: n7693_o = n7692_o;
      13'b0000000000001: n7693_o = n7692_o;
      default: n7693_o = n7692_o;
    endcase
  assign n7694_o = n1870_o[67];
  assign n7695_o = {n7694_o, n1978_o, n2137_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7696_o = n7695_o;
      13'b0100000000000: n7696_o = n7695_o;
      13'b0010000000000: n7696_o = n7695_o;
      13'b0001000000000: n7696_o = n7695_o;
      13'b0000100000000: n7696_o = n7695_o;
      13'b0000010000000: n7696_o = n7695_o;
      13'b0000001000000: n7696_o = n7695_o;
      13'b0000000100000: n7696_o = n7695_o;
      13'b0000000010000: n7696_o = n7695_o;
      13'b0000000001000: n7696_o = n7695_o;
      13'b0000000000100: n7696_o = n5782_o;
      13'b0000000000010: n7696_o = n7695_o;
      13'b0000000000001: n7696_o = n7695_o;
      default: n7696_o = n7695_o;
    endcase
  assign n7697_o = n1870_o[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7698_o = n7697_o;
      13'b0100000000000: n7698_o = n7697_o;
      13'b0010000000000: n7698_o = n7697_o;
      13'b0001000000000: n7698_o = n7697_o;
      13'b0000100000000: n7698_o = n7697_o;
      13'b0000010000000: n7698_o = n7697_o;
      13'b0000001000000: n7698_o = n7697_o;
      13'b0000000100000: n7698_o = n7697_o;
      13'b0000000010000: n7698_o = n7697_o;
      13'b0000000001000: n7698_o = n7697_o;
      13'b0000000000100: n7698_o = n5784_o;
      13'b0000000000010: n7698_o = n7697_o;
      13'b0000000000001: n7698_o = n7697_o;
      default: n7698_o = n7697_o;
    endcase
  assign n7699_o = n1870_o[71];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7700_o = n7699_o;
      13'b0100000000000: n7700_o = n7377_o;
      13'b0010000000000: n7700_o = n7699_o;
      13'b0001000000000: n7700_o = n7699_o;
      13'b0000100000000: n7700_o = n7699_o;
      13'b0000010000000: n7700_o = n7699_o;
      13'b0000001000000: n7700_o = n7699_o;
      13'b0000000100000: n7700_o = n7699_o;
      13'b0000000010000: n7700_o = n7699_o;
      13'b0000000001000: n7700_o = n7699_o;
      13'b0000000000100: n7700_o = n5786_o;
      13'b0000000000010: n7700_o = n7699_o;
      13'b0000000000001: n7700_o = n3075_o;
      default: n7700_o = n7699_o;
    endcase
  assign n7701_o = n5789_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7702_o = n2130_o;
      13'b0100000000000: n7702_o = n2130_o;
      13'b0010000000000: n7702_o = n2130_o;
      13'b0001000000000: n7702_o = n2130_o;
      13'b0000100000000: n7702_o = n2130_o;
      13'b0000010000000: n7702_o = n2130_o;
      13'b0000001000000: n7702_o = n2130_o;
      13'b0000000100000: n7702_o = n2130_o;
      13'b0000000010000: n7702_o = n6098_o;
      13'b0000000001000: n7702_o = n6029_o;
      13'b0000000000100: n7702_o = n7701_o;
      13'b0000000000010: n7702_o = n3266_o;
      13'b0000000000001: n7702_o = n3076_o;
      default: n7702_o = n2130_o;
    endcase
  assign n7703_o = n5789_o[1];
  assign n7704_o = n1870_o[74];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7705_o = n7704_o;
      13'b0100000000000: n7705_o = n7704_o;
      13'b0010000000000: n7705_o = n7704_o;
      13'b0001000000000: n7705_o = n7704_o;
      13'b0000100000000: n7705_o = n7704_o;
      13'b0000010000000: n7705_o = n7704_o;
      13'b0000001000000: n7705_o = n7704_o;
      13'b0000000100000: n7705_o = n7704_o;
      13'b0000000010000: n7705_o = n7704_o;
      13'b0000000001000: n7705_o = n7704_o;
      13'b0000000000100: n7705_o = n7703_o;
      13'b0000000000010: n7705_o = n7704_o;
      13'b0000000000001: n7705_o = n7704_o;
      default: n7705_o = n7704_o;
    endcase
  assign n7706_o = n1870_o[80];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7707_o = n7706_o;
      13'b0100000000000: n7707_o = n7706_o;
      13'b0010000000000: n7707_o = n7706_o;
      13'b0001000000000: n7707_o = n7706_o;
      13'b0000100000000: n7707_o = n7706_o;
      13'b0000010000000: n7707_o = n7706_o;
      13'b0000001000000: n7707_o = n6433_o;
      13'b0000000100000: n7707_o = n7706_o;
      13'b0000000010000: n7707_o = n7706_o;
      13'b0000000001000: n7707_o = n7706_o;
      13'b0000000000100: n7707_o = n7706_o;
      13'b0000000000010: n7707_o = n7706_o;
      13'b0000000000001: n7707_o = n7706_o;
      default: n7707_o = n7706_o;
    endcase
  assign n7708_o = n1870_o[82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7709_o = n7708_o;
      13'b0100000000000: n7709_o = n7708_o;
      13'b0010000000000: n7709_o = n7708_o;
      13'b0001000000000: n7709_o = n7708_o;
      13'b0000100000000: n7709_o = n7708_o;
      13'b0000010000000: n7709_o = n7708_o;
      13'b0000001000000: n7709_o = n7708_o;
      13'b0000000100000: n7709_o = n7708_o;
      13'b0000000010000: n7709_o = n7708_o;
      13'b0000000001000: n7709_o = n7708_o;
      13'b0000000000100: n7709_o = n7708_o;
      13'b0000000000010: n7709_o = n7708_o;
      13'b0000000000001: n7709_o = n3078_o;
      default: n7709_o = n7708_o;
    endcase
  assign n7710_o = n1870_o[84];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7711_o = n7710_o;
      13'b0100000000000: n7711_o = n7710_o;
      13'b0010000000000: n7711_o = n7710_o;
      13'b0001000000000: n7711_o = n7710_o;
      13'b0000100000000: n7711_o = n7710_o;
      13'b0000010000000: n7711_o = n7710_o;
      13'b0000001000000: n7711_o = n7710_o;
      13'b0000000100000: n7711_o = n7710_o;
      13'b0000000010000: n7711_o = n7710_o;
      13'b0000000001000: n7711_o = n7710_o;
      13'b0000000000100: n7711_o = n7710_o;
      13'b0000000000010: n7711_o = n7710_o;
      13'b0000000000001: n7711_o = n3080_o;
      default: n7711_o = n7710_o;
    endcase
  assign n7712_o = n1870_o[85];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7713_o = n7712_o;
      13'b0100000000000: n7713_o = n7712_o;
      13'b0010000000000: n7713_o = n7026_o;
      13'b0001000000000: n7713_o = n7712_o;
      13'b0000100000000: n7713_o = n7712_o;
      13'b0000010000000: n7713_o = n7712_o;
      13'b0000001000000: n7713_o = n7712_o;
      13'b0000000100000: n7713_o = n7712_o;
      13'b0000000010000: n7713_o = n7712_o;
      13'b0000000001000: n7713_o = n7712_o;
      13'b0000000000100: n7713_o = n7712_o;
      13'b0000000000010: n7713_o = n7712_o;
      13'b0000000000001: n7713_o = n7712_o;
      default: n7713_o = n7712_o;
    endcase
  assign n7714_o = n1870_o[86];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7715_o = n7714_o;
      13'b0100000000000: n7715_o = n7714_o;
      13'b0010000000000: n7715_o = n7714_o;
      13'b0001000000000: n7715_o = n7714_o;
      13'b0000100000000: n7715_o = n7714_o;
      13'b0000010000000: n7715_o = n7714_o;
      13'b0000001000000: n7715_o = n7714_o;
      13'b0000000100000: n7715_o = n7714_o;
      13'b0000000010000: n7715_o = n7714_o;
      13'b0000000001000: n7715_o = n7714_o;
      13'b0000000000100: n7715_o = n7714_o;
      13'b0000000000010: n7715_o = n7714_o;
      13'b0000000000001: n7715_o = n3082_o;
      default: n7715_o = n7714_o;
    endcase
  assign n7718_o = n1870_o[16:1];
  assign n7719_o = n1870_o[21];
  assign n7720_o = n1870_o[23];
  assign n7725_o = n1870_o[33:30];
  assign n7727_o = n1870_o[35];
  assign n7731_o = n1870_o[45];
  assign n7744_o = n1870_o[68];
  assign n7745_o = n1870_o[72];
  assign n7746_o = n1870_o[70];
  assign n7750_o = n1870_o[81];
  assign n7754_o = n6120_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7756_o = 1'b0;
      13'b0100000000000: n7756_o = 1'b0;
      13'b0010000000000: n7756_o = 1'b0;
      13'b0001000000000: n7756_o = 1'b0;
      13'b0000100000000: n7756_o = 1'b0;
      13'b0000010000000: n7756_o = 1'b0;
      13'b0000001000000: n7756_o = 1'b0;
      13'b0000000100000: n7756_o = n7754_o;
      13'b0000000010000: n7756_o = 1'b0;
      13'b0000000001000: n7756_o = 1'b0;
      13'b0000000000100: n7756_o = n5793_o;
      13'b0000000000010: n7756_o = n3299_o;
      13'b0000000000001: n7756_o = n3084_o;
      default: n7756_o = 1'b0;
    endcase
  assign n7757_o = n6120_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7759_o = 1'b0;
      13'b0100000000000: n7759_o = 1'b0;
      13'b0010000000000: n7759_o = 1'b0;
      13'b0001000000000: n7759_o = 1'b0;
      13'b0000100000000: n7759_o = 1'b0;
      13'b0000010000000: n7759_o = 1'b0;
      13'b0000001000000: n7759_o = 1'b0;
      13'b0000000100000: n7759_o = n7757_o;
      13'b0000000010000: n7759_o = 1'b0;
      13'b0000000001000: n7759_o = 1'b0;
      13'b0000000000100: n7759_o = 1'b0;
      13'b0000000000010: n7759_o = 1'b0;
      13'b0000000000001: n7759_o = 1'b0;
      default: n7759_o = 1'b0;
    endcase
  assign n7760_o = n5795_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7762_o = 1'b0;
      13'b0100000000000: n7762_o = 1'b0;
      13'b0010000000000: n7762_o = 1'b0;
      13'b0001000000000: n7762_o = 1'b0;
      13'b0000100000000: n7762_o = 1'b0;
      13'b0000010000000: n7762_o = 1'b0;
      13'b0000001000000: n7762_o = 1'b0;
      13'b0000000100000: n7762_o = 1'b0;
      13'b0000000010000: n7762_o = 1'b0;
      13'b0000000001000: n7762_o = 1'b0;
      13'b0000000000100: n7762_o = n7760_o;
      13'b0000000000010: n7762_o = 1'b0;
      13'b0000000000001: n7762_o = 1'b0;
      default: n7762_o = 1'b0;
    endcase
  assign n7763_o = n5795_o[1];
  assign n7764_o = n6031_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7766_o = 1'b0;
      13'b0100000000000: n7766_o = 1'b0;
      13'b0010000000000: n7766_o = n7028_o;
      13'b0001000000000: n7766_o = 1'b0;
      13'b0000100000000: n7766_o = 1'b0;
      13'b0000010000000: n7766_o = n6557_o;
      13'b0000001000000: n7766_o = n6435_o;
      13'b0000000100000: n7766_o = 1'b0;
      13'b0000000010000: n7766_o = 1'b0;
      13'b0000000001000: n7766_o = n7764_o;
      13'b0000000000100: n7766_o = n7763_o;
      13'b0000000000010: n7766_o = 1'b0;
      13'b0000000000001: n7766_o = n3086_o;
      default: n7766_o = 1'b0;
    endcase
  assign n7767_o = n6031_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7769_o = 1'b0;
      13'b0100000000000: n7769_o = 1'b0;
      13'b0010000000000: n7769_o = 1'b0;
      13'b0001000000000: n7769_o = 1'b0;
      13'b0000100000000: n7769_o = 1'b0;
      13'b0000010000000: n7769_o = 1'b0;
      13'b0000001000000: n7769_o = 1'b0;
      13'b0000000100000: n7769_o = 1'b0;
      13'b0000000010000: n7769_o = 1'b0;
      13'b0000000001000: n7769_o = n7767_o;
      13'b0000000000100: n7769_o = 1'b0;
      13'b0000000000010: n7769_o = 1'b0;
      13'b0000000000001: n7769_o = 1'b0;
      default: n7769_o = 1'b0;
    endcase
  assign n7770_o = n3088_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7772_o = 1'b0;
      13'b0100000000000: n7772_o = 1'b0;
      13'b0010000000000: n7772_o = 1'b0;
      13'b0001000000000: n7772_o = 1'b0;
      13'b0000100000000: n7772_o = 1'b0;
      13'b0000010000000: n7772_o = 1'b0;
      13'b0000001000000: n7772_o = n6437_o;
      13'b0000000100000: n7772_o = 1'b0;
      13'b0000000010000: n7772_o = 1'b0;
      13'b0000000001000: n7772_o = 1'b0;
      13'b0000000000100: n7772_o = 1'b0;
      13'b0000000000010: n7772_o = 1'b0;
      13'b0000000000001: n7772_o = n7770_o;
      default: n7772_o = 1'b0;
    endcase
  assign n7773_o = n3088_o[1];
  assign n7774_o = n5797_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7776_o = 1'b0;
      13'b0100000000000: n7776_o = 1'b0;
      13'b0010000000000: n7776_o = n7030_o;
      13'b0001000000000: n7776_o = 1'b0;
      13'b0000100000000: n7776_o = 1'b0;
      13'b0000010000000: n7776_o = 1'b0;
      13'b0000001000000: n7776_o = 1'b0;
      13'b0000000100000: n7776_o = 1'b0;
      13'b0000000010000: n7776_o = 1'b0;
      13'b0000000001000: n7776_o = 1'b0;
      13'b0000000000100: n7776_o = n7774_o;
      13'b0000000000010: n7776_o = 1'b0;
      13'b0000000000001: n7776_o = n7773_o;
      default: n7776_o = 1'b0;
    endcase
  assign n7777_o = n3088_o[2];
  assign n7778_o = n5797_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7780_o = 1'b0;
      13'b0100000000000: n7780_o = 1'b0;
      13'b0010000000000: n7780_o = 1'b0;
      13'b0001000000000: n7780_o = n6770_o;
      13'b0000100000000: n7780_o = 1'b0;
      13'b0000010000000: n7780_o = 1'b0;
      13'b0000001000000: n7780_o = 1'b0;
      13'b0000000100000: n7780_o = 1'b0;
      13'b0000000010000: n7780_o = 1'b0;
      13'b0000000001000: n7780_o = 1'b0;
      13'b0000000000100: n7780_o = n7778_o;
      13'b0000000000010: n7780_o = 1'b0;
      13'b0000000000001: n7780_o = n7777_o;
      default: n7780_o = 1'b0;
    endcase
  assign n7781_o = n3088_o[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7783_o = 1'b0;
      13'b0100000000000: n7783_o = 1'b0;
      13'b0010000000000: n7783_o = 1'b0;
      13'b0001000000000: n7783_o = n6772_o;
      13'b0000100000000: n7783_o = 1'b0;
      13'b0000010000000: n7783_o = 1'b0;
      13'b0000001000000: n7783_o = 1'b0;
      13'b0000000100000: n7783_o = 1'b0;
      13'b0000000010000: n7783_o = 1'b0;
      13'b0000000001000: n7783_o = 1'b0;
      13'b0000000000100: n7783_o = 1'b0;
      13'b0000000000010: n7783_o = 1'b0;
      13'b0000000000001: n7783_o = n7781_o;
      default: n7783_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7785_o = 1'b0;
      13'b0100000000000: n7785_o = 1'b0;
      13'b0010000000000: n7785_o = 1'b0;
      13'b0001000000000: n7785_o = n6774_o;
      13'b0000100000000: n7785_o = 1'b0;
      13'b0000010000000: n7785_o = 1'b0;
      13'b0000001000000: n7785_o = 1'b0;
      13'b0000000100000: n7785_o = 1'b0;
      13'b0000000010000: n7785_o = 1'b0;
      13'b0000000001000: n7785_o = 1'b0;
      13'b0000000000100: n7785_o = 1'b0;
      13'b0000000000010: n7785_o = 1'b0;
      13'b0000000000001: n7785_o = 1'b0;
      default: n7785_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7787_o = 1'b0;
      13'b0100000000000: n7787_o = 1'b0;
      13'b0010000000000: n7787_o = 1'b0;
      13'b0001000000000: n7787_o = 1'b0;
      13'b0000100000000: n7787_o = 1'b0;
      13'b0000010000000: n7787_o = 1'b0;
      13'b0000001000000: n7787_o = 1'b0;
      13'b0000000100000: n7787_o = 1'b0;
      13'b0000000010000: n7787_o = 1'b0;
      13'b0000000001000: n7787_o = 1'b0;
      13'b0000000000100: n7787_o = n5798_o;
      13'b0000000000010: n7787_o = 1'b0;
      13'b0000000000001: n7787_o = 1'b0;
      default: n7787_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7789_o = 1'b0;
      13'b0100000000000: n7789_o = 1'b0;
      13'b0010000000000: n7789_o = n7032_o;
      13'b0001000000000: n7789_o = 1'b0;
      13'b0000100000000: n7789_o = 1'b0;
      13'b0000010000000: n7789_o = 1'b0;
      13'b0000001000000: n7789_o = 1'b0;
      13'b0000000100000: n7789_o = 1'b0;
      13'b0000000010000: n7789_o = 1'b0;
      13'b0000000001000: n7789_o = 1'b0;
      13'b0000000000100: n7789_o = 1'b0;
      13'b0000000000010: n7789_o = 1'b0;
      13'b0000000000001: n7789_o = 1'b0;
      default: n7789_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7791_o = 1'b0;
      13'b0100000000000: n7791_o = 1'b0;
      13'b0010000000000: n7791_o = 1'b0;
      13'b0001000000000: n7791_o = 1'b0;
      13'b0000100000000: n7791_o = 1'b0;
      13'b0000010000000: n7791_o = 1'b0;
      13'b0000001000000: n7791_o = n6439_o;
      13'b0000000100000: n7791_o = 1'b0;
      13'b0000000010000: n7791_o = 1'b0;
      13'b0000000001000: n7791_o = 1'b0;
      13'b0000000000100: n7791_o = n5800_o;
      13'b0000000000010: n7791_o = 1'b0;
      13'b0000000000001: n7791_o = 1'b0;
      default: n7791_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7793_o = 1'b0;
      13'b0100000000000: n7793_o = 1'b0;
      13'b0010000000000: n7793_o = 1'b0;
      13'b0001000000000: n7793_o = 1'b0;
      13'b0000100000000: n7793_o = 1'b0;
      13'b0000010000000: n7793_o = 1'b0;
      13'b0000001000000: n7793_o = 1'b0;
      13'b0000000100000: n7793_o = 1'b0;
      13'b0000000010000: n7793_o = 1'b0;
      13'b0000000001000: n7793_o = 1'b0;
      13'b0000000000100: n7793_o = 1'b0;
      13'b0000000000010: n7793_o = 1'b0;
      13'b0000000000001: n7793_o = n3090_o;
      default: n7793_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7795_o = 1'b0;
      13'b0100000000000: n7795_o = 1'b0;
      13'b0010000000000: n7795_o = 1'b0;
      13'b0001000000000: n7795_o = 1'b0;
      13'b0000100000000: n7795_o = 1'b0;
      13'b0000010000000: n7795_o = 1'b0;
      13'b0000001000000: n7795_o = 1'b0;
      13'b0000000100000: n7795_o = 1'b0;
      13'b0000000010000: n7795_o = 1'b0;
      13'b0000000001000: n7795_o = 1'b0;
      13'b0000000000100: n7795_o = n5802_o;
      13'b0000000000010: n7795_o = 1'b0;
      13'b0000000000001: n7795_o = 1'b0;
      default: n7795_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7797_o = 1'b0;
      13'b0100000000000: n7797_o = 1'b0;
      13'b0010000000000: n7797_o = 1'b0;
      13'b0001000000000: n7797_o = 1'b0;
      13'b0000100000000: n7797_o = 1'b0;
      13'b0000010000000: n7797_o = 1'b0;
      13'b0000001000000: n7797_o = 1'b0;
      13'b0000000100000: n7797_o = 1'b0;
      13'b0000000010000: n7797_o = 1'b0;
      13'b0000000001000: n7797_o = n6033_o;
      13'b0000000000100: n7797_o = 1'b0;
      13'b0000000000010: n7797_o = 1'b0;
      13'b0000000000001: n7797_o = 1'b0;
      default: n7797_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7799_o = 1'b0;
      13'b0100000000000: n7799_o = 1'b0;
      13'b0010000000000: n7799_o = n7034_o;
      13'b0001000000000: n7799_o = 1'b0;
      13'b0000100000000: n7799_o = 1'b0;
      13'b0000010000000: n7799_o = 1'b0;
      13'b0000001000000: n7799_o = 1'b0;
      13'b0000000100000: n7799_o = 1'b0;
      13'b0000000010000: n7799_o = 1'b0;
      13'b0000000001000: n7799_o = 1'b0;
      13'b0000000000100: n7799_o = 1'b0;
      13'b0000000000010: n7799_o = 1'b0;
      13'b0000000000001: n7799_o = 1'b0;
      default: n7799_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7801_o = 1'b0;
      13'b0100000000000: n7801_o = n7379_o;
      13'b0010000000000: n7801_o = 1'b0;
      13'b0001000000000: n7801_o = n6776_o;
      13'b0000100000000: n7801_o = 1'b0;
      13'b0000010000000: n7801_o = 1'b0;
      13'b0000001000000: n7801_o = n6441_o;
      13'b0000000100000: n7801_o = 1'b0;
      13'b0000000010000: n7801_o = 1'b0;
      13'b0000000001000: n7801_o = n6035_o;
      13'b0000000000100: n7801_o = n5804_o;
      13'b0000000000010: n7801_o = 1'b0;
      13'b0000000000001: n7801_o = n3092_o;
      default: n7801_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7803_o = 1'b0;
      13'b0100000000000: n7803_o = 1'b0;
      13'b0010000000000: n7803_o = 1'b0;
      13'b0001000000000: n7803_o = 1'b0;
      13'b0000100000000: n7803_o = 1'b0;
      13'b0000010000000: n7803_o = 1'b0;
      13'b0000001000000: n7803_o = 1'b0;
      13'b0000000100000: n7803_o = 1'b0;
      13'b0000000010000: n7803_o = 1'b0;
      13'b0000000001000: n7803_o = 1'b0;
      13'b0000000000100: n7803_o = n5806_o;
      13'b0000000000010: n7803_o = 1'b0;
      13'b0000000000001: n7803_o = 1'b0;
      default: n7803_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7805_o = 1'b0;
      13'b0100000000000: n7805_o = 1'b0;
      13'b0010000000000: n7805_o = 1'b0;
      13'b0001000000000: n7805_o = 1'b0;
      13'b0000100000000: n7805_o = 1'b0;
      13'b0000010000000: n7805_o = 1'b0;
      13'b0000001000000: n7805_o = 1'b0;
      13'b0000000100000: n7805_o = 1'b0;
      13'b0000000010000: n7805_o = 1'b0;
      13'b0000000001000: n7805_o = 1'b0;
      13'b0000000000100: n7805_o = n5808_o;
      13'b0000000000010: n7805_o = 1'b0;
      13'b0000000000001: n7805_o = 1'b0;
      default: n7805_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7807_o = 1'b0;
      13'b0100000000000: n7807_o = 1'b0;
      13'b0010000000000: n7807_o = 1'b0;
      13'b0001000000000: n7807_o = 1'b0;
      13'b0000100000000: n7807_o = 1'b0;
      13'b0000010000000: n7807_o = 1'b0;
      13'b0000001000000: n7807_o = 1'b0;
      13'b0000000100000: n7807_o = 1'b0;
      13'b0000000010000: n7807_o = 1'b0;
      13'b0000000001000: n7807_o = 1'b0;
      13'b0000000000100: n7807_o = n5810_o;
      13'b0000000000010: n7807_o = 1'b0;
      13'b0000000000001: n7807_o = 1'b0;
      default: n7807_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7809_o = 2'b00;
      13'b0100000000000: n7809_o = 2'b00;
      13'b0010000000000: n7809_o = 2'b00;
      13'b0001000000000: n7809_o = 2'b00;
      13'b0000100000000: n7809_o = 2'b00;
      13'b0000010000000: n7809_o = 2'b00;
      13'b0000001000000: n7809_o = 2'b00;
      13'b0000000100000: n7809_o = 2'b00;
      13'b0000000010000: n7809_o = 2'b00;
      13'b0000000001000: n7809_o = 2'b00;
      13'b0000000000100: n7809_o = n5813_o;
      13'b0000000000010: n7809_o = 2'b00;
      13'b0000000000001: n7809_o = 2'b00;
      default: n7809_o = 2'b00;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7811_o = 1'b0;
      13'b0100000000000: n7811_o = n7380_o;
      13'b0010000000000: n7811_o = n7036_o;
      13'b0001000000000: n7811_o = 1'b0;
      13'b0000100000000: n7811_o = 1'b0;
      13'b0000010000000: n7811_o = n6559_o;
      13'b0000001000000: n7811_o = n6442_o;
      13'b0000000100000: n7811_o = n6122_o;
      13'b0000000010000: n7811_o = 1'b0;
      13'b0000000001000: n7811_o = n6036_o;
      13'b0000000000100: n7811_o = n5815_o;
      13'b0000000000010: n7811_o = n3301_o;
      13'b0000000000001: n7811_o = n3093_o;
      default: n7811_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7813_o = 1'b0;
      13'b0100000000000: n7813_o = 1'b0;
      13'b0010000000000: n7813_o = n7038_o;
      13'b0001000000000: n7813_o = 1'b0;
      13'b0000100000000: n7813_o = 1'b0;
      13'b0000010000000: n7813_o = 1'b0;
      13'b0000001000000: n7813_o = 1'b0;
      13'b0000000100000: n7813_o = 1'b0;
      13'b0000000010000: n7813_o = 1'b0;
      13'b0000000001000: n7813_o = 1'b0;
      13'b0000000000100: n7813_o = 1'b0;
      13'b0000000000010: n7813_o = 1'b0;
      13'b0000000000001: n7813_o = 1'b0;
      default: n7813_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7815_o = 2'b00;
      13'b0100000000000: n7815_o = n7382_o;
      13'b0010000000000: n7815_o = 2'b00;
      13'b0001000000000: n7815_o = 2'b00;
      13'b0000100000000: n7815_o = 2'b00;
      13'b0000010000000: n7815_o = 2'b00;
      13'b0000001000000: n7815_o = 2'b00;
      13'b0000000100000: n7815_o = 2'b00;
      13'b0000000010000: n7815_o = 2'b00;
      13'b0000000001000: n7815_o = 2'b00;
      13'b0000000000100: n7815_o = 2'b00;
      13'b0000000000010: n7815_o = 2'b00;
      13'b0000000000001: n7815_o = 2'b00;
      default: n7815_o = 2'b00;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7817_o = 2'b00;
      13'b0100000000000: n7817_o = 2'b00;
      13'b0010000000000: n7817_o = 2'b00;
      13'b0001000000000: n7817_o = 2'b00;
      13'b0000100000000: n7817_o = 2'b00;
      13'b0000010000000: n7817_o = 2'b00;
      13'b0000001000000: n7817_o = n6444_o;
      13'b0000000100000: n7817_o = 2'b00;
      13'b0000000010000: n7817_o = 2'b00;
      13'b0000000001000: n7817_o = 2'b00;
      13'b0000000000100: n7817_o = 2'b00;
      13'b0000000000010: n7817_o = 2'b00;
      13'b0000000000001: n7817_o = 2'b00;
      default: n7817_o = 2'b00;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7819_o = 1'b0;
      13'b0100000000000: n7819_o = n7383_o;
      13'b0010000000000: n7819_o = 1'b0;
      13'b0001000000000: n7819_o = 1'b0;
      13'b0000100000000: n7819_o = 1'b0;
      13'b0000010000000: n7819_o = 1'b0;
      13'b0000001000000: n7819_o = 1'b0;
      13'b0000000100000: n7819_o = 1'b0;
      13'b0000000010000: n7819_o = 1'b0;
      13'b0000000001000: n7819_o = 1'b0;
      13'b0000000000100: n7819_o = 1'b0;
      13'b0000000000010: n7819_o = 1'b0;
      13'b0000000000001: n7819_o = 1'b0;
      default: n7819_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7821_o = 1'b0;
      13'b0100000000000: n7821_o = 1'b0;
      13'b0010000000000: n7821_o = 1'b0;
      13'b0001000000000: n7821_o = 1'b0;
      13'b0000100000000: n7821_o = 1'b0;
      13'b0000010000000: n7821_o = 1'b0;
      13'b0000001000000: n7821_o = 1'b0;
      13'b0000000100000: n7821_o = 1'b0;
      13'b0000000010000: n7821_o = 1'b0;
      13'b0000000001000: n7821_o = 1'b0;
      13'b0000000000100: n7821_o = n5816_o;
      13'b0000000000010: n7821_o = 1'b0;
      13'b0000000000001: n7821_o = 1'b0;
      default: n7821_o = 1'b0;
    endcase
  assign n7833_o = n7822_o[9];
  assign n7841_o = n7822_o[19:17];
  assign n7845_o = n7822_o[27];
  assign n7847_o = n7822_o[29];
  assign n7852_o = n7822_o[66:35];
  assign n7854_o = n7822_o[74:68];
  assign n7857_o = n7822_o[80:79];
  assign n7858_o = n7822_o[87:82];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1640:17  */
  always @*
    case (n7528_o)
      13'b1000000000000: n7859_o = n2139_o;
      13'b0100000000000: n7859_o = n7384_o;
      13'b0010000000000: n7859_o = n2139_o;
      13'b0001000000000: n7859_o = n6777_o;
      13'b0000100000000: n7859_o = n2139_o;
      13'b0000010000000: n7859_o = n2139_o;
      13'b0000001000000: n7859_o = n6445_o;
      13'b0000000100000: n7859_o = n2139_o;
      13'b0000000010000: n7859_o = n6099_o;
      13'b0000000001000: n7859_o = n6037_o;
      13'b0000000000100: n7859_o = n5817_o;
      13'b0000000000010: n7859_o = n3268_o;
      13'b0000000000001: n7859_o = n3094_o;
      default: n7859_o = n2139_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:36  */
  assign n7860_o = set_exec[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:44  */
  assign n7861_o = ~n7860_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:60  */
  assign n7862_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:63  */
  assign n7863_o = ~n7862_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:77  */
  assign n7864_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:89  */
  assign n7866_o = n7864_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:68  */
  assign n7867_o = n7863_o | n7866_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3186:49  */
  assign n7868_o = n7861_o & n7867_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7870_o = n7892_o ? 1'b1 : n7811_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3189:34  */
  assign n7871_o = opcode[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3194:42  */
  assign n7873_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3194:33  */
  assign n7875_o = n7873_o ? 1'b1 : n7556_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3197:33  */
  assign n7877_o = setexecopc ? 1'b1 : n7574_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7879_o = n7885_o ? 1'b1 : n7543_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3189:25  */
  assign n7880_o = n7871_o ? n7556_o : n7875_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3189:25  */
  assign n7882_o = n7871_o ? n7559_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3189:25  */
  assign n7883_o = n7871_o ? n7574_o : n7877_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7884_o = n7891_o ? 1'b1 : n7801_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7885_o = build_logical & n7871_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7886_o = build_logical ? n7880_o : n7556_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7887_o = build_logical ? n7882_o : n7559_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7888_o = build_logical ? n7883_o : n7574_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7890_o = build_logical ? 1'b1 : n7612_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7891_o = build_logical & n7871_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3184:17  */
  assign n7892_o = build_logical & n7868_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:34  */
  assign n7895_o = opcode[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3211:50  */
  assign n7896_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3211:62  */
  assign n7898_o = n7896_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7900_o = n7931_o ? 1'b1 : n7673_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7904_o = n7922_o ? 2'b10 : n7533_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7906_o = n7927_o ? 1'b1 : n7568_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7907_o = n7929_o ? 1'b1 : n7641_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7908_o = n7930_o ? 1'b1 : n7665_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3210:33  */
  assign n7909_o = decodeopc & n7898_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7911_o = n7935_o ? 7'b0100001 : n7859_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7913_o = n7895_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7914_o = n7895_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7916_o = n7895_o ? n7888_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7917_o = n7895_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7918_o = n7895_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7919_o = n7895_o & n7909_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7920_o = n7895_o ? n7870_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3209:25  */
  assign n7921_o = n7895_o & decodeopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7922_o = build_bcd & n7913_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7924_o = build_bcd ? 1'b1 : n7879_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7926_o = build_bcd ? 1'b1 : n7887_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7927_o = build_bcd & n7914_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7928_o = build_bcd ? n7916_o : n7888_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7929_o = build_bcd & n7917_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7930_o = build_bcd & n7918_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7931_o = build_bcd & n7919_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7932_o = build_bcd ? 1'b1 : n7884_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7933_o = build_bcd ? 1'b1 : n7803_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7934_o = build_bcd ? n7920_o : n7870_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3204:17  */
  assign n7935_o = build_bcd & n7921_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3231:33  */
  assign n7936_o = ~trapd;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3229:17  */
  assign n7938_o = n7939_o ? 1'b1 : n7547_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3229:17  */
  assign n7939_o = set_z_error & n7936_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3229:17  */
  assign n7941_o = set_z_error ? 1'b1 : n7606_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3242:25  */
  assign n7943_o = clkena_lw ? trapmake : trapd;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3242:25  */
  assign n7944_o = clkena_lw ? next_micro_state : micro_state;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3240:17  */
  assign n7945_o = reset ? trapd : n7943_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3240:17  */
  assign n7947_o = reset ? 7'b0000010 : n7944_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3249:33  */
  assign n7953_o = micro_state == 7'b0000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3254:33  */
  assign n7956_o = micro_state == 7'b0000011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3259:33  */
  assign n7959_o = micro_state == 7'b0000100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:49  */
  assign n7960_o = brief[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:52  */
  assign n7961_o = ~n7960_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:57  */
  assign n7963_o = n7961_o | 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:82  */
  assign n7964_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:85  */
  assign n7965_o = ~n7964_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:90  */
  assign n7967_o = n7965_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:75  */
  assign n7968_o = n7963_o | n7967_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3272:57  */
  assign n7970_o = brief[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3274:59  */
  assign n7971_o = exec[22];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3274:49  */
  assign n7973_o = n7971_o ? 1'b1 : n2123_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3272:49  */
  assign n7975_o = n7970_o ? 1'b1 : n2116_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3272:49  */
  assign n7976_o = n7970_o ? n2123_o : n7973_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3277:57  */
  assign n7977_o = brief[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3277:60  */
  assign n7978_o = ~n7977_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3280:65  */
  assign n7979_o = brief[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3280:57  */
  assign n7981_o = n7979_o ? 1'b1 : n7702_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3277:49  */
  assign n7983_o = n7978_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3277:49  */
  assign n7984_o = n7978_o ? n7702_o : n7981_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7986_o = n7968_o ? 2'b01 : n7983_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7989_o = n7968_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7992_o = n7968_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7993_o = n7968_o ? n2116_o : n7975_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7994_o = n7968_o ? n2123_o : n7976_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7995_o = n7968_o ? 1'b1 : n7746_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7996_o = n7968_o ? n7702_o : n7984_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3265:41  */
  assign n7999_o = n7968_o ? 7'b0000110 : 7'b0001011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3264:33  */
  assign n8001_o = micro_state == 7'b0000101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3287:33  */
  assign n8004_o = micro_state == 7'b0000110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3295:49  */
  assign n8005_o = brief[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3295:41  */
  assign n8008_o = n8005_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:49  */
  assign n8009_o = brief[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:52  */
  assign n8010_o = ~n8009_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:66  */
  assign n8011_o = brief[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:69  */
  assign n8012_o = ~n8011_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:57  */
  assign n8013_o = n8010_o & n8012_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3301:57  */
  assign n8015_o = brief[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3301:69  */
  assign n8017_o = n8015_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3301:49  */
  assign n8020_o = n8017_o ? 7'b0000110 : 7'b0001100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:57  */
  assign n8021_o = brief[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:69  */
  assign n8023_o = n8021_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:49  */
  assign n8027_o = n8023_o ? n7904_o : 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:49  */
  assign n8030_o = n8023_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:49  */
  assign n8032_o = n8023_o ? 1'b1 : n7534_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:49  */
  assign n8033_o = n8023_o ? 1'b1 : n2129_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:49  */
  assign n8034_o = n8023_o ? n7702_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3307:49  */
  assign n8036_o = n8023_o ? n7911_o : 7'b0001101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:41  */
  assign n8038_o = n8013_o ? 2'b01 : n8027_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:41  */
  assign n8040_o = n8013_o ? 1'b0 : n8030_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:41  */
  assign n8041_o = n8013_o ? n7534_o : n8032_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:41  */
  assign n8042_o = n8013_o ? n2129_o : n8033_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:41  */
  assign n8043_o = n8013_o ? 1'b1 : n7746_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:41  */
  assign n8044_o = n8013_o ? n7702_o : n8034_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3298:41  */
  assign n8045_o = n8013_o ? n8020_o : n8036_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3294:33  */
  assign n8047_o = micro_state == 7'b0001011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3318:33  */
  assign n8050_o = micro_state == 7'b0001100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3328:49  */
  assign n8052_o = brief[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3328:52  */
  assign n8053_o = ~n8052_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3331:57  */
  assign n8054_o = brief[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3331:49  */
  assign n8056_o = n8054_o ? 1'b1 : n7702_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3328:41  */
  assign n8058_o = n8053_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3328:41  */
  assign n8059_o = n8053_o ? n7702_o : n8056_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3325:33  */
  assign n8061_o = micro_state == 7'b0001101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3338:49  */
  assign n8062_o = brief[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3338:41  */
  assign n8065_o = n8062_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:49  */
  assign n8066_o = brief[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:52  */
  assign n8067_o = ~n8066_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:66  */
  assign n8068_o = brief[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:57  */
  assign n8069_o = n8067_o & n8068_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:41  */
  assign n8073_o = n8069_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:41  */
  assign n8075_o = n8069_o ? n7534_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:41  */
  assign n8076_o = n8069_o ? n2129_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:41  */
  assign n8077_o = n8069_o ? 1'b1 : n7746_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3341:41  */
  assign n8079_o = n8069_o ? 7'b0000110 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3337:33  */
  assign n8081_o = micro_state == 7'b0001110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3351:33  */
  assign n8083_o = micro_state == 7'b0000111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:49  */
  assign n8084_o = brief[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:52  */
  assign n8085_o = ~n8084_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:57  */
  assign n8087_o = n8085_o | 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:82  */
  assign n8088_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:85  */
  assign n8089_o = ~n8088_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:90  */
  assign n8091_o = n8089_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:75  */
  assign n8092_o = n8087_o | n8091_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3364:57  */
  assign n8094_o = brief[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3364:49  */
  assign n8096_o = n8094_o ? 1'b1 : n2116_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3369:57  */
  assign n8097_o = brief[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3369:60  */
  assign n8098_o = ~n8097_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3372:65  */
  assign n8099_o = brief[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3372:57  */
  assign n8101_o = n8099_o ? 1'b1 : n7702_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3369:49  */
  assign n8103_o = n8098_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3369:49  */
  assign n8104_o = n8098_o ? n7702_o : n8101_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:41  */
  assign n8106_o = n8092_o ? 2'b01 : n8103_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:41  */
  assign n8109_o = n8092_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:41  */
  assign n8112_o = n8092_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:41  */
  assign n8113_o = n8092_o ? n2116_o : n8096_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:41  */
  assign n8114_o = n8092_o ? 1'b1 : n7746_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:41  */
  assign n8115_o = n8092_o ? n7702_o : n8104_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3357:41  */
  assign n8118_o = n8092_o ? 7'b0010100 : 7'b0001111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3356:33  */
  assign n8120_o = micro_state == 7'b0010011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3379:33  */
  assign n8123_o = micro_state == 7'b0010100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3388:49  */
  assign n8124_o = brief[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3388:41  */
  assign n8127_o = n8124_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:49  */
  assign n8128_o = brief[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:52  */
  assign n8129_o = ~n8128_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:66  */
  assign n8130_o = brief[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:69  */
  assign n8131_o = ~n8130_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:57  */
  assign n8132_o = n8129_o & n8131_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3394:57  */
  assign n8134_o = brief[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3394:69  */
  assign n8136_o = n8134_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3394:49  */
  assign n8139_o = n8136_o ? 7'b0010100 : 7'b0010000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3400:57  */
  assign n8140_o = brief[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3400:69  */
  assign n8142_o = n8140_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3400:49  */
  assign n8147_o = n8142_o ? 2'b11 : 2'b10;
  assign n8148_o = n7696_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3400:49  */
  assign n8149_o = n8142_o ? n8148_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3400:49  */
  assign n8150_o = n8142_o ? n7702_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3400:49  */
  assign n8153_o = n8142_o ? 7'b0000001 : 7'b0010001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:41  */
  assign n8155_o = n8132_o ? 2'b01 : n8147_o;
  assign n8156_o = n7696_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:41  */
  assign n8157_o = n8132_o ? n8156_o : n8149_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:41  */
  assign n8158_o = n8132_o ? 1'b1 : n7746_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:41  */
  assign n8159_o = n8132_o ? n7702_o : n8150_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3391:41  */
  assign n8160_o = n8132_o ? n8139_o : n8153_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3387:33  */
  assign n8162_o = micro_state == 7'b0001111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3411:33  */
  assign n8166_o = micro_state == 7'b0010000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3422:49  */
  assign n8169_o = brief[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3422:52  */
  assign n8170_o = ~n8169_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3425:57  */
  assign n8171_o = brief[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3425:49  */
  assign n8173_o = n8171_o ? 1'b1 : n7702_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3422:41  */
  assign n8175_o = n8170_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3422:41  */
  assign n8176_o = n8170_o ? n7702_o : n8173_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3418:33  */
  assign n8178_o = micro_state == 7'b0010001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3433:49  */
  assign n8180_o = brief[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3433:41  */
  assign n8183_o = n8180_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3436:49  */
  assign n8184_o = brief[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3436:52  */
  assign n8185_o = ~n8184_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3436:66  */
  assign n8186_o = brief[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3436:57  */
  assign n8187_o = n8185_o & n8186_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3436:41  */
  assign n8191_o = n8187_o ? 2'b01 : 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3436:41  */
  assign n8192_o = n8187_o ? 1'b1 : n7746_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3436:41  */
  assign n8195_o = n8187_o ? 7'b0010100 : 7'b0000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3431:33  */
  assign n8197_o = micro_state == 7'b0010010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3447:41  */
  assign n8199_o = exe_condition ? 1'b1 : n7529_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3447:41  */
  assign n8202_o = exe_condition ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3447:41  */
  assign n8204_o = exe_condition ? 7'b0000001 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3446:33  */
  assign n8206_o = micro_state == 7'b0010101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3453:33  */
  assign n8208_o = micro_state == 7'b0010110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3458:54  */
  assign n8209_o = ~long_start;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3458:41  */
  assign n8212_o = n8209_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3457:33  */
  assign n8215_o = micro_state == 7'b0010111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3467:33  */
  assign n8217_o = micro_state == 7'b0011000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3471:57  */
  assign n8218_o = ~exe_condition;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3473:57  */
  assign n8219_o = c_out[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3471:41  */
  assign n8221_o = n8227_o ? 1'b1 : n7529_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3473:49  */
  assign n8224_o = n8219_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3471:41  */
  assign n8226_o = n8233_o ? 7'b0000001 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3471:41  */
  assign n8227_o = n8218_o & n8219_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3471:41  */
  assign n8230_o = n8218_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3471:41  */
  assign n8232_o = n8218_o ? n8224_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3471:41  */
  assign n8233_o = n8218_o & n8219_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3470:33  */
  assign n8235_o = micro_state == 7'b0011001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3480:33  */
  assign n8241_o = micro_state == 7'b1000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3489:50  */
  assign n8242_o = sndopc[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3492:58  */
  assign n8243_o = opcode[10:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3492:71  */
  assign n8245_o = n8243_o == 2'b00;
  assign n8247_o = n1870_o[88];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3489:41  */
  assign n8248_o = n8255_o ? 1'b1 : n8247_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3489:41  */
  assign n8250_o = n8242_o ? 2'b10 : n7532_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3489:41  */
  assign n8253_o = n8242_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3489:41  */
  assign n8255_o = n8242_o & n8245_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3487:33  */
  assign n8260_o = micro_state == 7'b1000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3504:50  */
  assign n8262_o = sndopc[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3504:41  */
  assign n8264_o = n8262_o ? 2'b10 : n7532_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3504:41  */
  assign n8267_o = n8262_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3511:61  */
  assign n8271_o = exec[88];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3512:50  */
  assign n8272_o = sndopc[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3512:41  */
  assign n8274_o = n8272_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3512:41  */
  assign n8276_o = n8272_o ? 7'b1000100 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3501:33  */
  assign n8278_o = micro_state == 7'b1000011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3516:33  */
  assign n8280_o = micro_state == 7'b1000100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3520:49  */
  assign n8281_o = flags[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3520:41  */
  assign n8283_o = n8281_o ? 1'b1 : n7941_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3519:33  */
  assign n8285_o = micro_state == 7'b1000101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3525:33  */
  assign n8287_o = micro_state == 7'b0110111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:49  */
  assign n8288_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8295_o = n8288_o ? 2'b11 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8298_o = n8288_o ? 1'b0 : 1'b1;
  assign n8299_o = n1870_o[27];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8300_o = n8288_o ? n8299_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8301_o = n8288_o ? n7636_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8302_o = n8288_o ? 1'b1 : n7645_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8303_o = n8288_o ? 1'b1 : n1886_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8304_o = n8288_o ? n7713_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3530:41  */
  assign n8306_o = n8288_o ? 7'b0000001 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3528:33  */
  assign n8308_o = micro_state == 7'b0111000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3544:63  */
  assign n8309_o = sndopc[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3542:33  */
  assign n8312_o = micro_state == 7'b0111001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3547:33  */
  assign n8318_o = micro_state == 7'b0111010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3555:33  */
  assign n8321_o = micro_state == 7'b0111011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3560:49  */
  assign n8322_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3560:41  */
  assign n8324_o = n8322_o ? 1'b1 : n7715_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3559:33  */
  assign n8330_o = micro_state == 7'b0111100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3570:33  */
  assign n8333_o = micro_state == 7'b0111101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:49  */
  assign n8334_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3579:71  */
  assign n8336_o = sndopc[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8344_o = n8334_o ? 2'b11 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8347_o = n8334_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8349_o = n8334_o ? n8336_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8352_o = n8334_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8354_o = n8334_o ? 1'b1 : n7571_o;
  assign n8355_o = n1870_o[27];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8356_o = n8334_o ? n8355_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8357_o = n8334_o ? n7636_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8358_o = n8334_o ? 1'b1 : n7645_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8359_o = n8334_o ? 1'b1 : n2129_o;
  assign n8360_o = n7696_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8361_o = n8334_o ? n8360_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8362_o = n8334_o ? n7709_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8363_o = n8334_o ? n7713_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3575:41  */
  assign n8366_o = n8334_o ? 7'b0111111 : 7'b1000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3574:33  */
  assign n8368_o = micro_state == 7'b0111110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3592:33  */
  assign n8372_o = micro_state == 7'b0111111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3599:33  */
  assign n8376_o = micro_state == 7'b1000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:58  */
  assign n8377_o = last_data_read[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:71  */
  assign n8379_o = n8377_o != 16'b0000000000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3607:58  */
  assign n8380_o = opcode[5:3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3607:70  */
  assign n8382_o = n8380_o == 3'b100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3609:63  */
  assign n8384_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:41  */
  assign n8386_o = n8391_o ? 1'b1 : n7636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3607:49  */
  assign n8387_o = n8382_o & n8384_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:41  */
  assign n8388_o = n8392_o ? 1'b1 : n7686_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:41  */
  assign n8390_o = n8379_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:41  */
  assign n8391_o = n8379_o & n8387_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:41  */
  assign n8392_o = n8379_o & n8382_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3605:41  */
  assign n8394_o = n8379_o ? 7'b0011011 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3604:33  */
  assign n8396_o = micro_state == 7'b0011010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3616:53  */
  assign n8397_o = ~movem_run;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3622:58  */
  assign n8400_o = opcode[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3622:62  */
  assign n8401_o = ~n8400_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3622:49  */
  assign n8405_o = n8401_o ? 2'b11 : 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3622:49  */
  assign n8406_o = n8401_o ? 1'b1 : n7645_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3616:41  */
  assign n8408_o = n8397_o ? 2'b01 : n8405_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3616:41  */
  assign n8409_o = n8397_o ? n7645_o : n8406_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3616:41  */
  assign n8410_o = n8397_o ? n7686_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3616:41  */
  assign n8411_o = n8397_o ? n7698_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3616:41  */
  assign n8413_o = n8397_o ? n7911_o : 7'b0011011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3615:33  */
  assign n8415_o = micro_state == 7'b0011011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3631:50  */
  assign n8416_o = opcode[5:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3631:62  */
  assign n8418_o = n8416_o != 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3631:41  */
  assign n8420_o = n8418_o ? 1'b1 : n7534_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3630:33  */
  assign n8422_o = micro_state == 7'b0011101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3636:50  */
  assign n8423_o = opcode[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3636:62  */
  assign n8425_o = n8423_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3636:41  */
  assign n8427_o = n8425_o ? 1'b1 : n7900_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3635:33  */
  assign n8432_o = micro_state == 7'b0011110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3646:50  */
  assign n8433_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3646:63  */
  assign n8435_o = n8433_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3646:41  */
  assign n8437_o = n8435_o ? 1'b1 : n7900_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3651:50  */
  assign n8439_o = opcode[7:6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3651:63  */
  assign n8441_o = n8439_o == 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3651:41  */
  assign n8444_o = n8441_o ? 2'b00 : 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3645:33  */
  assign n8447_o = micro_state == 7'b0011111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3661:33  */
  assign n8449_o = micro_state == 7'b0100000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3665:50  */
  assign n8450_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3665:63  */
  assign n8452_o = n8450_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3665:41  */
  assign n8454_o = n8452_o ? 1'b1 : n7900_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3664:33  */
  assign n8457_o = micro_state == 7'b0100001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3675:50  */
  assign n8458_o = opcode[11:9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3675:63  */
  assign n8460_o = n8458_o == 3'b111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3675:41  */
  assign n8462_o = n8460_o ? 1'b1 : n7900_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3674:33  */
  assign n8465_o = micro_state == 7'b0100010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3684:33  */
  assign n8469_o = micro_state == 7'b0100011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3690:33  */
  assign n8472_o = micro_state == 7'b0100100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3694:33  */
  assign n8475_o = micro_state == 7'b0100101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3699:33  */
  assign n8478_o = micro_state == 7'b0100110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3703:33  */
  assign n8481_o = micro_state == 7'b0110010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3720:71  */
  assign n8484_o = trap_interrupt | trap_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3720:89  */
  assign n8485_o = n8484_o | trap_berr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3720:49  */
  assign n8487_o = n8485_o ? 1'b1 : n7938_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3714:41  */
  assign n8490_o = use_vbr_stackframe ? 2'b01 : 2'b10;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3714:41  */
  assign n8491_o = use_vbr_stackframe ? n7938_o : n8487_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3714:41  */
  assign n8492_o = use_vbr_stackframe ? 1'b1 : n1919_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3714:41  */
  assign n8495_o = use_vbr_stackframe ? 7'b0110100 : 7'b0110101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3710:33  */
  assign n8497_o = micro_state == 7'b0110011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3728:63  */
  assign n8498_o = trap_interrupt | trap_trace;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3728:41  */
  assign n8500_o = n8498_o ? 1'b1 : n7938_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3727:33  */
  assign n8503_o = micro_state == 7'b0110100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3742:41  */
  assign n8507_o = trap_berr ? 7'b1000110 : 7'b0110110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3736:33  */
  assign n8509_o = micro_state == 7'b0110101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3747:33  */
  assign n8513_o = micro_state == 7'b0110110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3754:33  */
  assign n8516_o = micro_state == 7'b1000110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3761:33  */
  assign n8519_o = micro_state == 7'b1000111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3768:33  */
  assign n8522_o = micro_state == 7'b1001000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3789:62  */
  assign n8525_o = ~use_vbr_stackframe;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3789:76  */
  assign n8526_o = opcode[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3789:67  */
  assign n8527_o = n8525_o | n8526_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3789:41  */
  assign n8530_o = n8527_o ? 1'b1 : n7727_o;
  assign n8531_o = n7691_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3789:41  */
  assign n8532_o = n8527_o ? 1'b1 : n8531_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3783:33  */
  assign n8534_o = micro_state == 7'b0101011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3797:77  */
  assign n8536_o = opcode[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3797:80  */
  assign n8537_o = ~n8536_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3797:67  */
  assign n8538_o = use_vbr_stackframe & n8537_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3797:41  */
  assign n8541_o = n8538_o ? 2'b10 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3797:41  */
  assign n8543_o = n8538_o ? 1'b1 : n7545_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3797:41  */
  assign n8544_o = n8538_o ? 1'b1 : n7659_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3797:41  */
  assign n8547_o = n8538_o ? 7'b0101101 : 7'b0000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3794:33  */
  assign n8549_o = micro_state == 7'b0101100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3810:33  */
  assign n8551_o = micro_state == 7'b0101101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3817:56  */
  assign n8552_o = last_data_in[15:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3817:70  */
  assign n8554_o = n8552_o == 4'b0010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3817:41  */
  assign n8558_o = n8554_o ? 2'b10 : 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3817:41  */
  assign n8560_o = n8554_o ? 2'b10 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3817:41  */
  assign n8562_o = n8554_o ? 1'b1 : n7545_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3817:41  */
  assign n8563_o = n8554_o ? 1'b1 : n7659_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3817:41  */
  assign n8566_o = n8554_o ? 7'b0101111 : 7'b0000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3815:33  */
  assign n8568_o = micro_state == 7'b0101110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3828:33  */
  assign n8570_o = micro_state == 7'b0101111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3832:33  */
  assign n8572_o = micro_state == 7'b0110000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3834:33  */
  assign n8575_o = micro_state == 7'b0110001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:50  */
  assign n8577_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:63  */
  assign n8579_o = n8577_o == 12'b000000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:79  */
  assign n8580_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:92  */
  assign n8582_o = n8580_o == 12'b000000000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:71  */
  assign n8583_o = n8579_o | n8582_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:108  */
  assign n8584_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:121  */
  assign n8586_o = n8584_o == 12'b100000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:100  */
  assign n8587_o = n8583_o | n8586_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:137  */
  assign n8588_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:150  */
  assign n8590_o = n8588_o == 12'b100000000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:129  */
  assign n8591_o = n8587_o | n8590_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:48  */
  assign n8592_o = cpu[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:66  */
  assign n8593_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:79  */
  assign n8595_o = n8593_o == 12'b000000000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:95  */
  assign n8596_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:108  */
  assign n8598_o = n8596_o == 12'b100000000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:87  */
  assign n8599_o = n8595_o | n8598_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:124  */
  assign n8600_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:137  */
  assign n8602_o = n8600_o == 12'b100000000011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:116  */
  assign n8603_o = n8599_o | n8602_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:153  */
  assign n8604_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:166  */
  assign n8606_o = n8604_o == 12'b100000000100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:145  */
  assign n8607_o = n8603_o | n8606_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3842:56  */
  assign n8608_o = n8592_o & n8607_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:159  */
  assign n8609_o = n8591_o | n8608_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3843:58  */
  assign n8610_o = opcode[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3843:61  */
  assign n8611_o = ~n8610_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:41  */
  assign n8613_o = n8618_o ? 1'b1 : n7636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:41  */
  assign n8615_o = n8609_o ? n7584_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:41  */
  assign n8617_o = n8609_o ? n7941_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3841:41  */
  assign n8618_o = n8609_o & n8611_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3838:33  */
  assign n8620_o = micro_state == 7'b1001001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3859:50  */
  assign n8624_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3859:41  */
  assign n8626_o = n8624_o ? 1'b1 : n7640_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3862:50  */
  assign n8627_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3862:53  */
  assign n8628_o = ~n8627_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3862:41  */
  assign n8631_o = n8628_o ? 2'b10 : 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3854:33  */
  assign n8633_o = micro_state == 7'b1001010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3869:50  */
  assign n8634_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3869:41  */
  assign n8637_o = n8634_o ? 1'b1 : n7643_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3869:41  */
  assign n8638_o = n8634_o ? 1'b1 : n7686_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3873:50  */
  assign n8639_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3873:53  */
  assign n8640_o = ~n8639_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3873:41  */
  assign n8643_o = n8640_o ? 2'b10 : 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3868:33  */
  assign n8645_o = micro_state == 7'b1001011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3880:50  */
  assign n8646_o = opcode[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3884:58  */
  assign n8650_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3884:61  */
  assign n8651_o = ~n8650_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3884:49  */
  assign n8654_o = n8651_o ? 2'b10 : 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3880:41  */
  assign n8656_o = n8646_o ? n7531_o : 2'b01;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3880:41  */
  assign n8657_o = n8646_o ? n8654_o : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3880:41  */
  assign n8658_o = n8646_o ? 1'b1 : n7643_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3880:41  */
  assign n8659_o = n8646_o ? 1'b1 : n7686_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3880:41  */
  assign n8660_o = n8646_o ? 1'b1 : n7745_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3880:41  */
  assign n8662_o = n8646_o ? 7'b1001101 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3879:33  */
  assign n8664_o = micro_state == 7'b1001100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3894:50  */
  assign n8665_o = opcode[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3894:53  */
  assign n8666_o = ~n8665_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3894:41  */
  assign n8669_o = n8666_o ? 2'b10 : 2'b11;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3893:33  */
  assign n8671_o = micro_state == 7'b1001101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3900:33  */
  assign n8673_o = micro_state == 7'b1001110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3904:50  */
  assign n8674_o = opcode[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3904:59  */
  assign n8676_o = n8674_o | 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3904:41  */
  assign n8679_o = n8676_o ? 6'b001110 : 6'b011110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3903:33  */
  assign n8681_o = micro_state == 7'b1010001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3913:51  */
  assign n8684_o = rot_cnt == 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3913:41  */
  assign n8687_o = n8684_o ? 7'b1010011 : 7'b1010010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3911:33  */
  assign n8689_o = micro_state == 7'b1010010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3920:50  */
  assign n8690_o = opcode[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3920:54  */
  assign n8691_o = ~n8690_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3920:41  */
  assign n8693_o = n8691_o ? 1'b1 : n7709_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:50  */
  assign n8695_o = opcode[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:54  */
  assign n8696_o = ~n8695_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:59  */
  assign n8698_o = n8696_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3928:58  */
  assign n8700_o = sndopc[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:41  */
  assign n8702_o = n8706_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:41  */
  assign n8704_o = n8712_o ? 7'b1010100 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:41  */
  assign n8706_o = n8698_o & n8700_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:41  */
  assign n8708_o = n8698_o ? 1'b1 : n7571_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:41  */
  assign n8709_o = n8698_o ? 1'b1 : n7636_o;
  assign n8710_o = n7696_o[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:41  */
  assign n8711_o = n8698_o ? 1'b1 : n8710_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3925:41  */
  assign n8712_o = n8698_o & n8700_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3919:33  */
  assign n8714_o = micro_state == 7'b1010011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3935:33  */
  assign n8719_o = micro_state == 7'b1010100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3941:33  */
  assign n8721_o = micro_state == 7'b1010101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:51  */
  assign n8722_o = op2out[31:16];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:65  */
  assign n8724_o = n8722_o == 16'b0000000000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:83  */
  assign n8725_o = opcode[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:74  */
  assign n8726_o = n8724_o | n8725_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:92  */
  assign n8728_o = n8726_o | 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:117  */
  assign n8729_o = op2out[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:130  */
  assign n8731_o = n8729_o == 16'b0000000000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:107  */
  assign n8732_o = n8728_o & n8731_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:41  */
  assign n8735_o = n8732_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3945:41  */
  assign n8737_o = n8732_o ? n7911_o : 7'b1010111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3944:33  */
  assign n8740_o = micro_state == 7'b1010110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3953:50  */
  assign n8741_o = opcode[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3953:59  */
  assign n8743_o = n8741_o | 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3953:41  */
  assign n8746_o = n8743_o ? 6'b001101 : 6'b011101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3952:33  */
  assign n8748_o = micro_state == 7'b1010111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3962:51  */
  assign n8751_o = rot_cnt == 6'b000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3962:41  */
  assign n8754_o = n8751_o ? 7'b1011001 : 7'b1011000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3960:33  */
  assign n8756_o = micro_state == 7'b1011000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3968:51  */
  assign n8757_o = ~z_error;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3968:70  */
  assign n8758_o = ~set_v_flag;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3968:56  */
  assign n8759_o = n8757_o & n8758_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3968:41  */
  assign n8761_o = n8759_o ? 1'b1 : n7636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3971:50  */
  assign n8762_o = opcode[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3971:54  */
  assign n8763_o = ~n8762_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3971:59  */
  assign n8765_o = n8763_o & 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3971:41  */
  assign n8768_o = n8765_o ? 2'b01 : n7904_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3971:41  */
  assign n8771_o = n8765_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3971:41  */
  assign n8772_o = n8765_o ? 1'b1 : n7744_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3971:41  */
  assign n8774_o = n8765_o ? 7'b1011010 : n7911_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3967:33  */
  assign n8777_o = micro_state == 7'b1011001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3980:48  */
  assign n8778_o = exec[34];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3980:41  */
  assign n8781_o = n8778_o ? 1'b1 : n7636_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3980:41  */
  assign n8782_o = n8778_o ? n7671_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3979:33  */
  assign n8785_o = micro_state == 7'b1011010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3989:50  */
  assign n8786_o = op2out[5:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3989:62  */
  assign n8788_o = n8786_o != 6'b000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3990:70  */
  assign n8789_o = op2out[5:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3989:41  */
  assign n8791_o = n8788_o ? n8789_o : n7577_o;
  assign n8792_o = n7822_o[23];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3989:41  */
  assign n8793_o = n8788_o ? n8792_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3988:33  */
  assign n8795_o = micro_state == 7'b1001111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3995:33  */
  assign n8797_o = micro_state == 7'b1010000;
  assign n8798_o = {n8797_o, n8795_o, n8785_o, n8777_o, n8756_o, n8748_o, n8740_o, n8721_o, n8719_o, n8714_o, n8689_o, n8681_o, n8673_o, n8671_o, n8664_o, n8645_o, n8633_o, n8620_o, n8575_o, n8572_o, n8570_o, n8568_o, n8551_o, n8549_o, n8534_o, n8522_o, n8519_o, n8516_o, n8513_o, n8509_o, n8503_o, n8497_o, n8481_o, n8478_o, n8475_o, n8472_o, n8469_o, n8465_o, n8457_o, n8449_o, n8447_o, n8432_o, n8422_o, n8415_o, n8396_o, n8376_o, n8372_o, n8368_o, n8333_o, n8330_o, n8321_o, n8318_o, n8312_o, n8308_o, n8287_o, n8285_o, n8280_o, n8278_o, n8260_o, n8241_o, n8235_o, n8217_o, n8215_o, n8208_o, n8206_o, n8197_o, n8178_o, n8166_o, n8162_o, n8123_o, n8120_o, n8083_o, n8081_o, n8061_o, n8050_o, n8047_o, n8004_o, n8001_o, n7959_o, n7956_o, n7953_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8801_o = 1'b1;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8801_o = n8221_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8801_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8801_o = n8199_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8801_o = n7529_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8801_o = n7529_o;
      default: n8801_o = n7529_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8814_o = n8656_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8814_o = n8558_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8814_o = 2'b01;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8814_o = 2'b01;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8814_o = 2'b01;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8814_o = 2'b01;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8814_o = n8490_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8814_o = 2'b10;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8814_o = n8444_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8814_o = n7531_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8814_o = n7531_o;
      default: n8814_o = n7531_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8815_o = n8264_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8815_o = n8250_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8815_o = n7532_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8815_o = n7532_o;
      default: n8815_o = n7532_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n8768_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b01;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n8702_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n8669_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8853_o = n8657_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8853_o = n8643_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8853_o = n8631_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8853_o = n8560_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8853_o = n8541_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8853_o = n8408_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8853_o = n8390_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8853_o = n8344_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8853_o = n8295_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8853_o = n8274_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8853_o = 2'b01;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8853_o = n8191_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8853_o = n8175_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8853_o = 2'b10;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8853_o = n8155_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8853_o = n8106_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8853_o = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8853_o = n8073_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8853_o = n8058_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8853_o = 2'b10;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8853_o = n8038_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8853_o = n7986_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8853_o = n7904_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8853_o = 2'b11;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8853_o = n7904_o;
      default: n8853_o = n7904_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8856_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8856_o = n8040_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8856_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8856_o = 1'b0;
      default: n8856_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8859_o = n8230_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8859_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8859_o = 1'b0;
      default: n8859_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8864_o = n8420_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8864_o = n8075_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8864_o = n8041_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8864_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8864_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8864_o = n7534_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8864_o = 1'b1;
      default: n8864_o = n7534_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8866_o = n8109_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8866_o = n7989_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8866_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8866_o = 1'b0;
      default: n8866_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8876_o = n8183_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8876_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8876_o = n8127_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8876_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8876_o = n8112_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8876_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8876_o = n8065_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8876_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8876_o = n8008_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8876_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8876_o = n7992_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8876_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8876_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8876_o = 1'b0;
      default: n8876_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8880_o = n8232_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8880_o = n8212_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8880_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8880_o = n8202_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8880_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8880_o = 1'b0;
      default: n8880_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8894_o = n8562_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8894_o = n8543_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8894_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8894_o = n7545_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8894_o = n7545_o;
      default: n8894_o = n7545_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8896_o = n8500_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8896_o = n8491_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8896_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8896_o = n7938_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8896_o = n7938_o;
      default: n8896_o = n7938_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b1;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8899_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8899_o = 1'b0;
      default: n8899_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8902_o = 1'b1;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8902_o = n7886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8902_o = n7886_o;
      default: n8902_o = n7886_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8905_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8905_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8905_o = 1'b0;
      default: n8905_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8909_o = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8909_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8909_o = 1'b0;
      default: n8909_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8913_o = n8347_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8913_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8913_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8913_o = 1'b0;
      default: n8913_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8916_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8916_o = n7565_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8916_o = n7565_o;
      default: n8916_o = n7565_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8921_o = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8921_o = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8921_o = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8921_o = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8921_o = n7906_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8921_o = n7906_o;
      default: n8921_o = n7906_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8923_o = n8349_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8923_o = n8309_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8923_o = n8267_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8923_o = n8253_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8923_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8923_o = 1'b0;
      default: n8923_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8928_o = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8928_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8928_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8928_o = 1'b0;
      default: n8928_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8931_o = n8352_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8931_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8931_o = 1'b0;
      default: n8931_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = 1'b1;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n8708_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8937_o = n8354_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8937_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8937_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8937_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8937_o = n7571_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8937_o = n7571_o;
      default: n8937_o = n7571_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = n8771_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8941_o = 1'b1;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8941_o = n8298_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8941_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8941_o = 1'b0;
      default: n8941_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8946_o = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8946_o = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8946_o = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8946_o = n7928_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8946_o = n7928_o;
      default: n8946_o = n7928_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n8791_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n8746_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n8679_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8947_o = n7577_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8947_o = n7577_o;
      default: n8947_o = n7577_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8951_o = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8951_o = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8951_o = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8951_o = n7581_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8951_o = n7581_o;
      default: n8951_o = n7581_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8954_o = 1'b1;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8954_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8954_o = 1'b0;
      default: n8954_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8961_o = 1'b1;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8961_o = 1'b1;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8961_o = 1'b1;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8961_o = 1'b1;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8961_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8961_o = 1'b0;
      default: n8961_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8963_o = n8615_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8963_o = n7584_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8963_o = n7584_o;
      default: n8963_o = n7584_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8964_o = n8617_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8964_o = n8283_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8964_o = n7941_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8964_o = n7941_o;
      default: n8964_o = n7941_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8967_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8967_o = n8113_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8967_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8967_o = n7993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8967_o = n2116_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8967_o = n2116_o;
      default: n8967_o = n2116_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = n8735_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8969_o = 1'b0;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8969_o = 1'b0;
      default: n8969_o = 1'b0;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8971_o = 1'b1;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8971_o = n7624_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8971_o = n7624_o;
      default: n8971_o = n7624_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = 1'b1;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8972_o = n7628_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8972_o = n7628_o;
      default: n8972_o = n7628_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = 1'b1;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = 1'b1;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8973_o = n7719_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8973_o = n7719_o;
      default: n8973_o = n7719_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8974_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8974_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8974_o = n7994_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8974_o = n2123_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8974_o = n2123_o;
      default: n8974_o = n2123_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = 1'b1;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8975_o = n7630_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8975_o = n7630_o;
      default: n8975_o = n7630_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8976_o = n8492_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8976_o = n1919_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8976_o = n1919_o;
      default: n8976_o = n1919_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8977_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8977_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8977_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8977_o = n7632_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8977_o = n7632_o;
      default: n8977_o = n7632_o;
    endcase
  assign n8978_o = n1870_o[27];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8979_o = 1'b1;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8979_o = 1'b1;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8979_o = n8356_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8979_o = n8300_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8979_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8979_o = n8978_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8979_o = n8978_o;
      default: n8979_o = n8978_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n8781_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n8761_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n8709_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8980_o = n8613_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8980_o = 1'b1;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8980_o = 1'b1;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8980_o = n8386_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8980_o = 1'b1;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8980_o = n8357_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8980_o = n8301_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8980_o = n7636_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8980_o = n7636_o;
      default: n8980_o = n7636_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8981_o = 1'b1;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8981_o = n8530_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8981_o = n7727_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8981_o = n7727_o;
      default: n8981_o = n7727_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8982_o = n8626_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8982_o = n7640_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8982_o = n7640_o;
      default: n8982_o = n7640_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8983_o = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8983_o = n7907_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8983_o = n7907_o;
      default: n8983_o = n7907_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8984_o = n8658_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8984_o = n8637_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8984_o = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8984_o = n7643_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8984_o = n7643_o;
      default: n8984_o = n7643_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8985_o = n8409_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8985_o = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8985_o = n8358_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8985_o = n8302_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8985_o = n7645_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8985_o = n7645_o;
      default: n8985_o = n7645_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8986_o = n7731_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8986_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8986_o = 1'b1;
      default: n8986_o = n7731_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8987_o = n8563_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8987_o = n8544_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8987_o = 1'b1;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8987_o = 1'b1;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8987_o = 1'b1;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8987_o = n7659_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8987_o = n7659_o;
      default: n8987_o = n7659_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8988_o = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8988_o = n7908_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8988_o = n7908_o;
      default: n8988_o = n7908_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n8782_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8989_o = n7671_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8989_o = n7671_o;
      default: n8989_o = n7671_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8990_o = n8462_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8990_o = n8454_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8990_o = n8437_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8990_o = n8427_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8990_o = n7900_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8990_o = n7900_o;
      default: n8990_o = n7900_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8991_o = n8659_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8991_o = n8638_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8991_o = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8991_o = n8410_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8991_o = n8388_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8991_o = n7686_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8991_o = n7686_o;
      default: n8991_o = n7686_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8992_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8992_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8992_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8992_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8992_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8992_o = n7689_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8992_o = n7689_o;
      default: n8992_o = n7689_o;
    endcase
  assign n8993_o = n7691_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8994_o = 1'b1;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8994_o = 1'b1;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8994_o = n8993_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8994_o = n8993_o;
      default: n8994_o = n8993_o;
    endcase
  assign n8995_o = n7691_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8996_o = n8532_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8996_o = 1'b1;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8996_o = n8995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8996_o = n8995_o;
      default: n8996_o = n8995_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8997_o = 1'b1;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8997_o = n8359_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8997_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8997_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8997_o = n8076_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8997_o = n8042_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8997_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8997_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8997_o = n2129_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8997_o = 1'b1;
      default: n8997_o = n2129_o;
    endcase
  assign n8998_o = n7696_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8999_o = n8361_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8999_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8999_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8999_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8999_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8999_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8999_o = n8157_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8999_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8999_o = n8998_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8999_o = n8998_o;
      default: n8999_o = n8998_o;
    endcase
  assign n9000_o = n7696_o[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n8711_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9001_o = n9000_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9001_o = n9000_o;
      default: n9001_o = n9000_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n8772_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = 1'b1;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9002_o = n7744_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9002_o = n7744_o;
      default: n9002_o = n7744_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9003_o = n8411_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9003_o = n7698_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9003_o = n7698_o;
      default: n9003_o = n7698_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9004_o = 1'b1;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9004_o = n8192_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9004_o = n8158_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9004_o = n8114_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9004_o = n8077_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9004_o = n8043_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9004_o = n7995_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9004_o = n7746_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9004_o = n7746_o;
      default: n9004_o = n7746_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9005_o = n8660_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9005_o = 1'b1;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9005_o = n7745_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9005_o = n7745_o;
      default: n9005_o = n7745_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9006_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9006_o = n8176_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9006_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9006_o = n8159_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9006_o = n8115_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9006_o = n8059_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9006_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9006_o = n8044_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9006_o = n7996_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9006_o = n7702_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9006_o = n7702_o;
      default: n9006_o = n7702_o;
    endcase
  assign n9007_o = n1870_o[79];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9008_o = 1'b1;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9008_o = 1'b1;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9008_o = n9007_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9008_o = n9007_o;
      default: n9008_o = n9007_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n8693_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9009_o = n8362_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9009_o = n7709_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9009_o = n7709_o;
      default: n9009_o = n7709_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9010_o = n8303_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9010_o = n1886_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9010_o = n1886_o;
      default: n9010_o = n1886_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9011_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9011_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9011_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9011_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9011_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9011_o = n7711_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9011_o = n7711_o;
      default: n9011_o = n7711_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9012_o = 1'b1;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9012_o = n8363_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9012_o = n8304_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9012_o = n7713_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9012_o = n7713_o;
      default: n9012_o = n7713_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9013_o = n8324_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9013_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9013_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9013_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9013_o = n7715_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9013_o = n7715_o;
      default: n9013_o = n7715_o;
    endcase
  assign n9014_o = n1870_o[87];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9015_o = 1'b1;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9015_o = n9014_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9015_o = n9014_o;
      default: n9015_o = n9014_o;
    endcase
  assign n9016_o = n1870_o[88];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9017_o = n8271_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9017_o = n8248_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9017_o = n9016_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9017_o = n9016_o;
      default: n9017_o = n9016_o;
    endcase
  assign n9018_o = n1870_o[28];
  assign n9020_o = n7691_o[3:2];
  assign n9022_o = n7696_o[0];
  assign n9023_o = n7696_o[3:2];
  assign n9024_o = n1870_o[78:75];
  assign n9026_o = n7822_o[23];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n8793_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9027_o = n9026_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9027_o = n9026_o;
      default: n9027_o = n9026_o;
    endcase
  assign n9028_o = n7822_o[25:24];
  assign n9029_o = n7822_o[22:21];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3248:25  */
  always @*
    case (n8798_o)
      81'b100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n8774_o;
      81'b000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n8754_o;
      81'b000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b1011000;
      81'b000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n8737_o;
      81'b000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b1010110;
      81'b000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n8704_o;
      81'b000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n8687_o;
      81'b000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b1010010;
      81'b000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b1001110;
      81'b000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9070_o = n8662_o;
      81'b000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b1001100;
      81'b000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b1001011;
      81'b000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b0110001;
      81'b000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b0000001;
      81'b000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9070_o = n8566_o;
      81'b000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9070_o = 7'b0101110;
      81'b000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9070_o = n8547_o;
      81'b000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9070_o = 7'b0101100;
      81'b000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9070_o = 7'b0110110;
      81'b000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9070_o = 7'b1001000;
      81'b000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9070_o = 7'b1000111;
      81'b000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9070_o = 7'b0011000;
      81'b000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9070_o = n8507_o;
      81'b000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9070_o = 7'b0110101;
      81'b000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9070_o = n8495_o;
      81'b000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9070_o = 7'b0110011;
      81'b000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9070_o = 7'b0100110;
      81'b000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9070_o = 7'b0100100;
      81'b000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9070_o = 7'b0100000;
      81'b000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9070_o = 7'b0011111;
      81'b000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9070_o = n8413_o;
      81'b000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9070_o = n8394_o;
      81'b000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9070_o = 7'b0011000;
      81'b000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9070_o = n8366_o;
      81'b000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9070_o = 7'b0111110;
      81'b000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9070_o = 7'b0111101;
      81'b000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9070_o = 7'b0111100;
      81'b000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9070_o = 7'b0111011;
      81'b000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9070_o = 7'b0111010;
      81'b000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9070_o = n8306_o;
      81'b000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9070_o = 7'b0111000;
      81'b000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9070_o = 7'b1000101;
      81'b000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9070_o = n8276_o;
      81'b000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9070_o = 7'b1000011;
      81'b000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9070_o = 7'b1000010;
      81'b000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9070_o = n8226_o;
      81'b000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9070_o = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9070_o = 7'b0011000;
      81'b000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9070_o = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9070_o = n8204_o;
      81'b000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9070_o = n8195_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9070_o = 7'b0010010;
      81'b000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9070_o = 7'b0010001;
      81'b000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9070_o = n8160_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9070_o = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9070_o = n8118_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9070_o = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9070_o = n8079_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9070_o = 7'b0001110;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9070_o = 7'b0001101;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9070_o = n8045_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9070_o = n7999_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9070_o = n7911_o;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9070_o = 7'b0000001;
      81'b000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9070_o = n7911_o;
      default: n9070_o = n7911_o;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4012:41  */
  assign n9076_o = exec[33];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4012:33  */
  assign n9077_o = clkena_lw & n9076_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4013:27  */
  assign n9078_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4014:47  */
  assign n9079_o = reg_qa[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4014:19  */
  assign n9081_o = n9078_o == 12'b000000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4015:47  */
  assign n9082_o = reg_qa[2:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4015:19  */
  assign n9084_o = n9078_o == 12'b000000000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4016:48  */
  assign n9085_o = reg_qa[3:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4016:19  */
  assign n9087_o = n9078_o == 12'b000000000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4017:19  */
  assign n9089_o = n9078_o == 12'b100000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4018:19  */
  assign n9091_o = n9078_o == 12'b100000000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4019:19  */
  assign n9093_o = n9078_o == 12'b100000000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4020:19  */
  assign n9095_o = n9078_o == 12'b100000000011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4021:19  */
  assign n9097_o = n9078_o == 12'b100000000100;
  assign n9098_o = {n9097_o, n9095_o, n9093_o, n9091_o, n9089_o, n9087_o, n9084_o, n9081_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n9098_o)
      8'b10000000: n9099_o = vbr;
      8'b01000000: n9099_o = vbr;
      8'b00100000: n9099_o = vbr;
      8'b00010000: n9099_o = reg_qa;
      8'b00001000: n9099_o = vbr;
      8'b00000100: n9099_o = vbr;
      8'b00000010: n9099_o = vbr;
      8'b00000001: n9099_o = vbr;
      default: n9099_o = vbr;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n9098_o)
      8'b10000000: n9100_o = cacr;
      8'b01000000: n9100_o = cacr;
      8'b00100000: n9100_o = cacr;
      8'b00010000: n9100_o = cacr;
      8'b00001000: n9100_o = cacr;
      8'b00000100: n9100_o = n9085_o;
      8'b00000010: n9100_o = cacr;
      8'b00000001: n9100_o = cacr;
      default: n9100_o = cacr;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n9098_o)
      8'b10000000: n9101_o = dfc;
      8'b01000000: n9101_o = dfc;
      8'b00100000: n9101_o = dfc;
      8'b00010000: n9101_o = dfc;
      8'b00001000: n9101_o = dfc;
      8'b00000100: n9101_o = dfc;
      8'b00000010: n9101_o = n9082_o;
      8'b00000001: n9101_o = dfc;
      default: n9101_o = dfc;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4013:17  */
  always @*
    case (n9098_o)
      8'b10000000: n9102_o = sfc;
      8'b01000000: n9102_o = sfc;
      8'b00100000: n9102_o = sfc;
      8'b00010000: n9102_o = sfc;
      8'b00001000: n9102_o = sfc;
      8'b00000100: n9102_o = sfc;
      8'b00000010: n9102_o = sfc;
      8'b00000001: n9102_o = n9079_o;
      default: n9102_o = sfc;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4012:11  */
  assign n9103_o = n9077_o ? n9099_o : vbr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4012:11  */
  assign n9104_o = n9077_o ? n9100_o : cacr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4012:11  */
  assign n9105_o = n9077_o ? n9101_o : dfc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4012:11  */
  assign n9106_o = n9077_o ? n9102_o : sfc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4009:11  */
  assign n9108_o = reset ? 32'b00000000000000000000000000000000 : n9103_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4009:11  */
  assign n9110_o = reset ? 4'b0000 : n9104_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4009:11  */
  assign n9111_o = reset ? dfc : n9105_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4009:11  */
  assign n9112_o = reset ? sfc : n9106_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4028:19  */
  assign n9117_o = brief[11:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4029:78  */
  assign n9119_o = {29'b00000000000000000000000000000, sfc};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4029:17  */
  assign n9121_o = n9117_o == 12'b000000000000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4030:78  */
  assign n9123_o = {29'b00000000000000000000000000000, dfc};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4030:17  */
  assign n9125_o = n9117_o == 12'b000000000001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4031:79  */
  assign n9127_o = cacr & 4'b0011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4031:71  */
  assign n9129_o = {28'b0000000000000000000000000000, n9127_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4031:11  */
  assign n9131_o = n9117_o == 12'b000000000010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4033:11  */
  assign n9133_o = n9117_o == 12'b100000000001;
  assign n9134_o = {n9133_o, n9131_o, n9125_o, n9121_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4028:9  */
  always @*
    case (n9134_o)
      4'b1000: n9136_o = vbr;
      4'b0100: n9136_o = n9129_o;
      4'b0010: n9136_o = n9123_o;
      4'b0001: n9136_o = n9119_o;
      default: n9136_o = 32'b00000000000000000000000000000000;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4047:32  */
  assign n9141_o = exe_opcode[11:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4048:25  */
  assign n9143_o = n9141_o == 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4049:25  */
  assign n9145_o = n9141_o == 4'b0001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4050:65  */
  assign n9146_o = flags[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4050:56  */
  assign n9147_o = ~n9146_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4050:82  */
  assign n9148_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4050:73  */
  assign n9149_o = ~n9148_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4050:69  */
  assign n9150_o = n9147_o & n9149_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4050:25  */
  assign n9152_o = n9141_o == 4'b0010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4051:60  */
  assign n9153_o = flags[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4051:72  */
  assign n9154_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4051:64  */
  assign n9155_o = n9153_o | n9154_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4051:25  */
  assign n9157_o = n9141_o == 4'b0011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4052:64  */
  assign n9158_o = flags[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4052:55  */
  assign n9159_o = ~n9158_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4052:25  */
  assign n9161_o = n9141_o == 4'b0100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4053:60  */
  assign n9162_o = flags[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4053:25  */
  assign n9164_o = n9141_o == 4'b0101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4054:64  */
  assign n9165_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4054:55  */
  assign n9166_o = ~n9165_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4054:25  */
  assign n9168_o = n9141_o == 4'b0110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4055:60  */
  assign n9169_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4055:25  */
  assign n9171_o = n9141_o == 4'b0111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4056:64  */
  assign n9172_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4056:55  */
  assign n9173_o = ~n9172_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4056:25  */
  assign n9175_o = n9141_o == 4'b1000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4057:60  */
  assign n9176_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4057:25  */
  assign n9178_o = n9141_o == 4'b1001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4058:64  */
  assign n9179_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4058:55  */
  assign n9180_o = ~n9179_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4058:25  */
  assign n9182_o = n9141_o == 4'b1010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4059:60  */
  assign n9183_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4059:25  */
  assign n9185_o = n9141_o == 4'b1011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:61  */
  assign n9186_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:74  */
  assign n9187_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:65  */
  assign n9188_o = n9186_o & n9187_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:92  */
  assign n9189_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:83  */
  assign n9190_o = ~n9189_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:109  */
  assign n9191_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:100  */
  assign n9192_o = ~n9191_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:96  */
  assign n9193_o = n9190_o & n9192_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:79  */
  assign n9194_o = n9188_o | n9193_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4060:25  */
  assign n9196_o = n9141_o == 4'b1100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:61  */
  assign n9197_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:78  */
  assign n9198_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:69  */
  assign n9199_o = ~n9198_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:65  */
  assign n9200_o = n9197_o & n9199_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:96  */
  assign n9201_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:87  */
  assign n9202_o = ~n9201_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:109  */
  assign n9203_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:100  */
  assign n9204_o = n9202_o & n9203_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:83  */
  assign n9205_o = n9200_o | n9204_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4061:25  */
  assign n9207_o = n9141_o == 4'b1101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:61  */
  assign n9208_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:74  */
  assign n9209_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:65  */
  assign n9210_o = n9208_o & n9209_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:91  */
  assign n9211_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:82  */
  assign n9212_o = ~n9211_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:78  */
  assign n9213_o = n9210_o & n9212_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:109  */
  assign n9214_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:100  */
  assign n9215_o = ~n9214_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:126  */
  assign n9216_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:117  */
  assign n9217_o = ~n9216_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:113  */
  assign n9218_o = n9215_o & n9217_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:143  */
  assign n9219_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:134  */
  assign n9220_o = ~n9219_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:130  */
  assign n9221_o = n9218_o & n9220_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:96  */
  assign n9222_o = n9213_o | n9221_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4062:25  */
  assign n9224_o = n9141_o == 4'b1110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:61  */
  assign n9225_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:78  */
  assign n9226_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:69  */
  assign n9227_o = ~n9226_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:65  */
  assign n9228_o = n9225_o & n9227_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:96  */
  assign n9229_o = flags[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:87  */
  assign n9230_o = ~n9229_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:109  */
  assign n9231_o = flags[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:100  */
  assign n9232_o = n9230_o & n9231_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:83  */
  assign n9233_o = n9228_o | n9232_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:122  */
  assign n9234_o = flags[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:114  */
  assign n9235_o = n9233_o | n9234_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4063:25  */
  assign n9237_o = n9141_o == 4'b1111;
  assign n9238_o = {n9237_o, n9224_o, n9207_o, n9196_o, n9185_o, n9182_o, n9178_o, n9175_o, n9171_o, n9168_o, n9164_o, n9161_o, n9157_o, n9152_o, n9145_o, n9143_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4047:17  */
  always @*
    case (n9238_o)
      16'b1000000000000000: n9241_o = n9235_o;
      16'b0100000000000000: n9241_o = n9222_o;
      16'b0010000000000000: n9241_o = n9205_o;
      16'b0001000000000000: n9241_o = n9194_o;
      16'b0000100000000000: n9241_o = n9183_o;
      16'b0000010000000000: n9241_o = n9180_o;
      16'b0000001000000000: n9241_o = n9176_o;
      16'b0000000100000000: n9241_o = n9173_o;
      16'b0000000010000000: n9241_o = n9169_o;
      16'b0000000001000000: n9241_o = n9166_o;
      16'b0000000000100000: n9241_o = n9162_o;
      16'b0000000000010000: n9241_o = n9159_o;
      16'b0000000000001000: n9241_o = n9155_o;
      16'b0000000000000100: n9241_o = n9150_o;
      16'b0000000000000010: n9241_o = 1'b0;
      16'b0000000000000001: n9241_o = 1'b1;
      default: n9241_o = exe_condition;
    endcase
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4075:54  */
  assign n9246_o = exec[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4077:60  */
  assign n9247_o = data_read[15:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4078:43  */
  assign n9248_o = exec[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4078:68  */
  assign n9249_o = set[69];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4078:62  */
  assign n9250_o = n9248_o | n9249_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4080:49  */
  assign n9253_o = movem_regaddr == 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4081:49  */
  assign n9256_o = movem_regaddr == 4'b0001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4082:49  */
  assign n9259_o = movem_regaddr == 4'b0010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4083:49  */
  assign n9262_o = movem_regaddr == 4'b0011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4084:49  */
  assign n9265_o = movem_regaddr == 4'b0100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4085:49  */
  assign n9268_o = movem_regaddr == 4'b0101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4086:49  */
  assign n9271_o = movem_regaddr == 4'b0110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4087:49  */
  assign n9274_o = movem_regaddr == 4'b0111;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4088:49  */
  assign n9277_o = movem_regaddr == 4'b1000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4089:49  */
  assign n9280_o = movem_regaddr == 4'b1001;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4090:49  */
  assign n9283_o = movem_regaddr == 4'b1010;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4091:49  */
  assign n9286_o = movem_regaddr == 4'b1011;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4092:49  */
  assign n9289_o = movem_regaddr == 4'b1100;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4093:49  */
  assign n9292_o = movem_regaddr == 4'b1101;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4094:49  */
  assign n9295_o = movem_regaddr == 4'b1110;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4095:49  */
  assign n9298_o = movem_regaddr == 4'b1111;
  assign n9299_o = {n9298_o, n9295_o, n9292_o, n9289_o, n9286_o, n9283_o, n9280_o, n9277_o, n9274_o, n9271_o, n9268_o, n9265_o, n9262_o, n9259_o, n9256_o, n9253_o};
  assign n9300_o = sndopc[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9301_o = n9300_o;
      16'b0100000000000000: n9301_o = n9300_o;
      16'b0010000000000000: n9301_o = n9300_o;
      16'b0001000000000000: n9301_o = n9300_o;
      16'b0000100000000000: n9301_o = n9300_o;
      16'b0000010000000000: n9301_o = n9300_o;
      16'b0000001000000000: n9301_o = n9300_o;
      16'b0000000100000000: n9301_o = n9300_o;
      16'b0000000010000000: n9301_o = n9300_o;
      16'b0000000001000000: n9301_o = n9300_o;
      16'b0000000000100000: n9301_o = n9300_o;
      16'b0000000000010000: n9301_o = n9300_o;
      16'b0000000000001000: n9301_o = n9300_o;
      16'b0000000000000100: n9301_o = n9300_o;
      16'b0000000000000010: n9301_o = n9300_o;
      16'b0000000000000001: n9301_o = 1'b0;
      default: n9301_o = n9300_o;
    endcase
  assign n9302_o = sndopc[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9303_o = n9302_o;
      16'b0100000000000000: n9303_o = n9302_o;
      16'b0010000000000000: n9303_o = n9302_o;
      16'b0001000000000000: n9303_o = n9302_o;
      16'b0000100000000000: n9303_o = n9302_o;
      16'b0000010000000000: n9303_o = n9302_o;
      16'b0000001000000000: n9303_o = n9302_o;
      16'b0000000100000000: n9303_o = n9302_o;
      16'b0000000010000000: n9303_o = n9302_o;
      16'b0000000001000000: n9303_o = n9302_o;
      16'b0000000000100000: n9303_o = n9302_o;
      16'b0000000000010000: n9303_o = n9302_o;
      16'b0000000000001000: n9303_o = n9302_o;
      16'b0000000000000100: n9303_o = n9302_o;
      16'b0000000000000010: n9303_o = 1'b0;
      16'b0000000000000001: n9303_o = n9302_o;
      default: n9303_o = n9302_o;
    endcase
  assign n9304_o = sndopc[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9305_o = n9304_o;
      16'b0100000000000000: n9305_o = n9304_o;
      16'b0010000000000000: n9305_o = n9304_o;
      16'b0001000000000000: n9305_o = n9304_o;
      16'b0000100000000000: n9305_o = n9304_o;
      16'b0000010000000000: n9305_o = n9304_o;
      16'b0000001000000000: n9305_o = n9304_o;
      16'b0000000100000000: n9305_o = n9304_o;
      16'b0000000010000000: n9305_o = n9304_o;
      16'b0000000001000000: n9305_o = n9304_o;
      16'b0000000000100000: n9305_o = n9304_o;
      16'b0000000000010000: n9305_o = n9304_o;
      16'b0000000000001000: n9305_o = n9304_o;
      16'b0000000000000100: n9305_o = 1'b0;
      16'b0000000000000010: n9305_o = n9304_o;
      16'b0000000000000001: n9305_o = n9304_o;
      default: n9305_o = n9304_o;
    endcase
  assign n9306_o = sndopc[3];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9307_o = n9306_o;
      16'b0100000000000000: n9307_o = n9306_o;
      16'b0010000000000000: n9307_o = n9306_o;
      16'b0001000000000000: n9307_o = n9306_o;
      16'b0000100000000000: n9307_o = n9306_o;
      16'b0000010000000000: n9307_o = n9306_o;
      16'b0000001000000000: n9307_o = n9306_o;
      16'b0000000100000000: n9307_o = n9306_o;
      16'b0000000010000000: n9307_o = n9306_o;
      16'b0000000001000000: n9307_o = n9306_o;
      16'b0000000000100000: n9307_o = n9306_o;
      16'b0000000000010000: n9307_o = n9306_o;
      16'b0000000000001000: n9307_o = 1'b0;
      16'b0000000000000100: n9307_o = n9306_o;
      16'b0000000000000010: n9307_o = n9306_o;
      16'b0000000000000001: n9307_o = n9306_o;
      default: n9307_o = n9306_o;
    endcase
  assign n9308_o = sndopc[4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9309_o = n9308_o;
      16'b0100000000000000: n9309_o = n9308_o;
      16'b0010000000000000: n9309_o = n9308_o;
      16'b0001000000000000: n9309_o = n9308_o;
      16'b0000100000000000: n9309_o = n9308_o;
      16'b0000010000000000: n9309_o = n9308_o;
      16'b0000001000000000: n9309_o = n9308_o;
      16'b0000000100000000: n9309_o = n9308_o;
      16'b0000000010000000: n9309_o = n9308_o;
      16'b0000000001000000: n9309_o = n9308_o;
      16'b0000000000100000: n9309_o = n9308_o;
      16'b0000000000010000: n9309_o = 1'b0;
      16'b0000000000001000: n9309_o = n9308_o;
      16'b0000000000000100: n9309_o = n9308_o;
      16'b0000000000000010: n9309_o = n9308_o;
      16'b0000000000000001: n9309_o = n9308_o;
      default: n9309_o = n9308_o;
    endcase
  assign n9310_o = sndopc[5];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9311_o = n9310_o;
      16'b0100000000000000: n9311_o = n9310_o;
      16'b0010000000000000: n9311_o = n9310_o;
      16'b0001000000000000: n9311_o = n9310_o;
      16'b0000100000000000: n9311_o = n9310_o;
      16'b0000010000000000: n9311_o = n9310_o;
      16'b0000001000000000: n9311_o = n9310_o;
      16'b0000000100000000: n9311_o = n9310_o;
      16'b0000000010000000: n9311_o = n9310_o;
      16'b0000000001000000: n9311_o = n9310_o;
      16'b0000000000100000: n9311_o = 1'b0;
      16'b0000000000010000: n9311_o = n9310_o;
      16'b0000000000001000: n9311_o = n9310_o;
      16'b0000000000000100: n9311_o = n9310_o;
      16'b0000000000000010: n9311_o = n9310_o;
      16'b0000000000000001: n9311_o = n9310_o;
      default: n9311_o = n9310_o;
    endcase
  assign n9312_o = sndopc[6];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9313_o = n9312_o;
      16'b0100000000000000: n9313_o = n9312_o;
      16'b0010000000000000: n9313_o = n9312_o;
      16'b0001000000000000: n9313_o = n9312_o;
      16'b0000100000000000: n9313_o = n9312_o;
      16'b0000010000000000: n9313_o = n9312_o;
      16'b0000001000000000: n9313_o = n9312_o;
      16'b0000000100000000: n9313_o = n9312_o;
      16'b0000000010000000: n9313_o = n9312_o;
      16'b0000000001000000: n9313_o = 1'b0;
      16'b0000000000100000: n9313_o = n9312_o;
      16'b0000000000010000: n9313_o = n9312_o;
      16'b0000000000001000: n9313_o = n9312_o;
      16'b0000000000000100: n9313_o = n9312_o;
      16'b0000000000000010: n9313_o = n9312_o;
      16'b0000000000000001: n9313_o = n9312_o;
      default: n9313_o = n9312_o;
    endcase
  assign n9314_o = sndopc[7];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9315_o = n9314_o;
      16'b0100000000000000: n9315_o = n9314_o;
      16'b0010000000000000: n9315_o = n9314_o;
      16'b0001000000000000: n9315_o = n9314_o;
      16'b0000100000000000: n9315_o = n9314_o;
      16'b0000010000000000: n9315_o = n9314_o;
      16'b0000001000000000: n9315_o = n9314_o;
      16'b0000000100000000: n9315_o = n9314_o;
      16'b0000000010000000: n9315_o = 1'b0;
      16'b0000000001000000: n9315_o = n9314_o;
      16'b0000000000100000: n9315_o = n9314_o;
      16'b0000000000010000: n9315_o = n9314_o;
      16'b0000000000001000: n9315_o = n9314_o;
      16'b0000000000000100: n9315_o = n9314_o;
      16'b0000000000000010: n9315_o = n9314_o;
      16'b0000000000000001: n9315_o = n9314_o;
      default: n9315_o = n9314_o;
    endcase
  assign n9316_o = sndopc[8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9317_o = n9316_o;
      16'b0100000000000000: n9317_o = n9316_o;
      16'b0010000000000000: n9317_o = n9316_o;
      16'b0001000000000000: n9317_o = n9316_o;
      16'b0000100000000000: n9317_o = n9316_o;
      16'b0000010000000000: n9317_o = n9316_o;
      16'b0000001000000000: n9317_o = n9316_o;
      16'b0000000100000000: n9317_o = 1'b0;
      16'b0000000010000000: n9317_o = n9316_o;
      16'b0000000001000000: n9317_o = n9316_o;
      16'b0000000000100000: n9317_o = n9316_o;
      16'b0000000000010000: n9317_o = n9316_o;
      16'b0000000000001000: n9317_o = n9316_o;
      16'b0000000000000100: n9317_o = n9316_o;
      16'b0000000000000010: n9317_o = n9316_o;
      16'b0000000000000001: n9317_o = n9316_o;
      default: n9317_o = n9316_o;
    endcase
  assign n9318_o = sndopc[9];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9319_o = n9318_o;
      16'b0100000000000000: n9319_o = n9318_o;
      16'b0010000000000000: n9319_o = n9318_o;
      16'b0001000000000000: n9319_o = n9318_o;
      16'b0000100000000000: n9319_o = n9318_o;
      16'b0000010000000000: n9319_o = n9318_o;
      16'b0000001000000000: n9319_o = 1'b0;
      16'b0000000100000000: n9319_o = n9318_o;
      16'b0000000010000000: n9319_o = n9318_o;
      16'b0000000001000000: n9319_o = n9318_o;
      16'b0000000000100000: n9319_o = n9318_o;
      16'b0000000000010000: n9319_o = n9318_o;
      16'b0000000000001000: n9319_o = n9318_o;
      16'b0000000000000100: n9319_o = n9318_o;
      16'b0000000000000010: n9319_o = n9318_o;
      16'b0000000000000001: n9319_o = n9318_o;
      default: n9319_o = n9318_o;
    endcase
  assign n9320_o = sndopc[10];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9321_o = n9320_o;
      16'b0100000000000000: n9321_o = n9320_o;
      16'b0010000000000000: n9321_o = n9320_o;
      16'b0001000000000000: n9321_o = n9320_o;
      16'b0000100000000000: n9321_o = n9320_o;
      16'b0000010000000000: n9321_o = 1'b0;
      16'b0000001000000000: n9321_o = n9320_o;
      16'b0000000100000000: n9321_o = n9320_o;
      16'b0000000010000000: n9321_o = n9320_o;
      16'b0000000001000000: n9321_o = n9320_o;
      16'b0000000000100000: n9321_o = n9320_o;
      16'b0000000000010000: n9321_o = n9320_o;
      16'b0000000000001000: n9321_o = n9320_o;
      16'b0000000000000100: n9321_o = n9320_o;
      16'b0000000000000010: n9321_o = n9320_o;
      16'b0000000000000001: n9321_o = n9320_o;
      default: n9321_o = n9320_o;
    endcase
  assign n9322_o = sndopc[11];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9323_o = n9322_o;
      16'b0100000000000000: n9323_o = n9322_o;
      16'b0010000000000000: n9323_o = n9322_o;
      16'b0001000000000000: n9323_o = n9322_o;
      16'b0000100000000000: n9323_o = 1'b0;
      16'b0000010000000000: n9323_o = n9322_o;
      16'b0000001000000000: n9323_o = n9322_o;
      16'b0000000100000000: n9323_o = n9322_o;
      16'b0000000010000000: n9323_o = n9322_o;
      16'b0000000001000000: n9323_o = n9322_o;
      16'b0000000000100000: n9323_o = n9322_o;
      16'b0000000000010000: n9323_o = n9322_o;
      16'b0000000000001000: n9323_o = n9322_o;
      16'b0000000000000100: n9323_o = n9322_o;
      16'b0000000000000010: n9323_o = n9322_o;
      16'b0000000000000001: n9323_o = n9322_o;
      default: n9323_o = n9322_o;
    endcase
  assign n9324_o = sndopc[12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9325_o = n9324_o;
      16'b0100000000000000: n9325_o = n9324_o;
      16'b0010000000000000: n9325_o = n9324_o;
      16'b0001000000000000: n9325_o = 1'b0;
      16'b0000100000000000: n9325_o = n9324_o;
      16'b0000010000000000: n9325_o = n9324_o;
      16'b0000001000000000: n9325_o = n9324_o;
      16'b0000000100000000: n9325_o = n9324_o;
      16'b0000000010000000: n9325_o = n9324_o;
      16'b0000000001000000: n9325_o = n9324_o;
      16'b0000000000100000: n9325_o = n9324_o;
      16'b0000000000010000: n9325_o = n9324_o;
      16'b0000000000001000: n9325_o = n9324_o;
      16'b0000000000000100: n9325_o = n9324_o;
      16'b0000000000000010: n9325_o = n9324_o;
      16'b0000000000000001: n9325_o = n9324_o;
      default: n9325_o = n9324_o;
    endcase
  assign n9326_o = sndopc[13];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9327_o = n9326_o;
      16'b0100000000000000: n9327_o = n9326_o;
      16'b0010000000000000: n9327_o = 1'b0;
      16'b0001000000000000: n9327_o = n9326_o;
      16'b0000100000000000: n9327_o = n9326_o;
      16'b0000010000000000: n9327_o = n9326_o;
      16'b0000001000000000: n9327_o = n9326_o;
      16'b0000000100000000: n9327_o = n9326_o;
      16'b0000000010000000: n9327_o = n9326_o;
      16'b0000000001000000: n9327_o = n9326_o;
      16'b0000000000100000: n9327_o = n9326_o;
      16'b0000000000010000: n9327_o = n9326_o;
      16'b0000000000001000: n9327_o = n9326_o;
      16'b0000000000000100: n9327_o = n9326_o;
      16'b0000000000000010: n9327_o = n9326_o;
      16'b0000000000000001: n9327_o = n9326_o;
      default: n9327_o = n9326_o;
    endcase
  assign n9328_o = sndopc[14];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9329_o = n9328_o;
      16'b0100000000000000: n9329_o = 1'b0;
      16'b0010000000000000: n9329_o = n9328_o;
      16'b0001000000000000: n9329_o = n9328_o;
      16'b0000100000000000: n9329_o = n9328_o;
      16'b0000010000000000: n9329_o = n9328_o;
      16'b0000001000000000: n9329_o = n9328_o;
      16'b0000000100000000: n9329_o = n9328_o;
      16'b0000000010000000: n9329_o = n9328_o;
      16'b0000000001000000: n9329_o = n9328_o;
      16'b0000000000100000: n9329_o = n9328_o;
      16'b0000000000010000: n9329_o = n9328_o;
      16'b0000000000001000: n9329_o = n9328_o;
      16'b0000000000000100: n9329_o = n9328_o;
      16'b0000000000000010: n9329_o = n9328_o;
      16'b0000000000000001: n9329_o = n9328_o;
      default: n9329_o = n9328_o;
    endcase
  assign n9330_o = sndopc[15];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4079:41  */
  always @*
    case (n9299_o)
      16'b1000000000000000: n9331_o = 1'b0;
      16'b0100000000000000: n9331_o = n9330_o;
      16'b0010000000000000: n9331_o = n9330_o;
      16'b0001000000000000: n9331_o = n9330_o;
      16'b0000100000000000: n9331_o = n9330_o;
      16'b0000010000000000: n9331_o = n9330_o;
      16'b0000001000000000: n9331_o = n9330_o;
      16'b0000000100000000: n9331_o = n9330_o;
      16'b0000000010000000: n9331_o = n9330_o;
      16'b0000000001000000: n9331_o = n9330_o;
      16'b0000000000100000: n9331_o = n9330_o;
      16'b0000000000010000: n9331_o = n9330_o;
      16'b0000000000001000: n9331_o = n9330_o;
      16'b0000000000000100: n9331_o = n9330_o;
      16'b0000000000000010: n9331_o = n9330_o;
      16'b0000000000000001: n9331_o = n9330_o;
      default: n9331_o = n9330_o;
    endcase
  assign n9332_o = {n9331_o, n9329_o, n9327_o, n9325_o, n9323_o, n9321_o, n9319_o, n9317_o, n9315_o, n9313_o, n9311_o, n9309_o, n9307_o, n9305_o, n9303_o, n9301_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4078:33  */
  assign n9333_o = n9250_o ? n9332_o : sndopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4076:33  */
  assign n9334_o = decodeopc ? n9247_o : n9333_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4107:26  */
  assign n9342_o = sndopc[3:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4107:38  */
  assign n9344_o = n9342_o == 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4108:34  */
  assign n9345_o = sndopc[7:4];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4108:46  */
  assign n9347_o = n9345_o == 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4110:42  */
  assign n9349_o = sndopc[11:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4110:55  */
  assign n9351_o = n9349_o == 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4111:50  */
  assign n9352_o = sndopc[15:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4111:64  */
  assign n9354_o = n9352_o == 4'b0000;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4111:41  */
  assign n9357_o = n9354_o ? 1'b0 : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4115:60  */
  assign n9359_o = sndopc[15:12];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4117:60  */
  assign n9360_o = sndopc[11:8];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4110:33  */
  assign n9362_o = n9351_o ? 1'b1 : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4110:33  */
  assign n9363_o = n9351_o ? n9359_o : n9360_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4110:33  */
  assign n9365_o = n9351_o ? n9357_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4120:52  */
  assign n9366_o = sndopc[7:4];
  assign n9368_o = {1'b1, n9362_o};
  assign n9369_o = n9368_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4108:25  */
  assign n9370_o = n9347_o ? n9369_o : 1'b1;
  assign n9371_o = n9368_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4108:25  */
  assign n9373_o = n9347_o ? n9371_o : 1'b0;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4108:25  */
  assign n9374_o = n9347_o ? n9363_o : n9366_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4108:25  */
  assign n9376_o = n9347_o ? n9365_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4124:44  */
  assign n9377_o = sndopc[3:0];
  assign n9378_o = {n9373_o, n9370_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4107:17  */
  assign n9380_o = n9344_o ? n9378_o : 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4107:17  */
  assign n9383_o = n9344_o ? n9374_o : n9377_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4107:17  */
  assign n9385_o = n9344_o ? n9376_o : 1'b1;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4126:29  */
  assign n9387_o = movem_mux[1:0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4126:41  */
  assign n9389_o = n9387_o == 2'b00;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4128:37  */
  assign n9391_o = movem_mux[2];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4128:40  */
  assign n9392_o = ~n9391_o;
  assign n9394_o = n9381_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4128:25  */
  assign n9395_o = n9392_o ? 1'b1 : n9394_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4132:37  */
  assign n9396_o = movem_mux[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4132:40  */
  assign n9397_o = ~n9396_o;
  assign n9399_o = n9381_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4132:25  */
  assign n9400_o = n9397_o ? 1'b1 : n9399_o;
  assign n9401_o = {1'b1, n9395_o};
  assign n9402_o = n9401_o[0];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4126:17  */
  assign n9403_o = n9389_o ? n9402_o : n9400_o;
  assign n9404_o = n9401_o[1];
  assign n9405_o = n9381_o[1];
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4126:17  */
  assign n9406_o = n9389_o ? n9404_o : n9405_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:464:17  */
  always @(posedge clk)
    n9409_q <= n106_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:458:17  */
  assign n9410_o = clkena_in ? n87_o : syncreset;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n83_o)
    if (n83_o)
      n9411_q <= 4'b0000;
    else
      n9411_q <= n9410_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:458:17  */
  assign n9412_o = clkena_in ? n89_o : reset;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n83_o)
    if (n83_o)
      n9413_q <= 1'b1;
    else
      n9413_q <= n9412_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9414_q <= n1473_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  assign n9415_o = n1023_o ? addr : tmp_tg68_pc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9416_q <= n9415_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  assign n9417_o = n1024_o ? addr : memaddr;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9418_q <= n9417_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9419_q <= n1475_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9420_q <= n1476_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9421_q <= n1478_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9422_q <= n1480_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9423_q <= n1481_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4073:17  */
  assign n9424_o = clkena_lw ? n9334_o : sndopc;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4073:17  */
  always @(posedge clk)
    n9425_q <= n9424_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9426_q <= n1482_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9427_q <= n1483_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9428_q <= n1485_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  assign n9430_o = clkena_lw ? rf_source_addr : rf_source_addrd;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9431_q <= n9430_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  assign n9432_o = {n337_o, n316_o, n334_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  assign n9435_o = clkena_lw ? rf_dest_addr : rdindex_a;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9436_q <= n9435_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  assign n9437_o = clkena_lw ? rf_source_addr : rdindex_b;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9438_q <= n9437_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  assign n9439_o = clkena_lw ? n272_o : wr_areg;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9440_q <= n9439_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  assign n9441_o = clkena_in ? n1010_o : memaddr_delta_rega;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9442_q <= n9441_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  assign n9443_o = clkena_in ? n1012_o : memaddr_delta_regb;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9444_q <= n9443_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  assign n9445_o = clkena_in ? n1015_o : use_base;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:941:17  */
  always @(posedge clk)
    n9446_q <= n9445_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9447_q <= n751_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  assign n9448_o = {n600_o, n607_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9450_q <= n752_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9451_q <= n1486_o;
  assign n9453_o = {n948_o, n945_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9454_q <= n1488_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9455_q <= n1489_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9456_q <= n754_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9457_q <= n1491_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9458_q <= n1493_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9459_q <= n756_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9460_q <= n1495_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9461_q <= n1497_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9462_q <= n1499_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9463_q <= n1845_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9464_q <= n757_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1254:17  */
  assign n9465_o = clkena_lw ? n1608_o : exec_tas;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1254:17  */
  always @(posedge clk)
    n9466_q <= n9465_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9467_q <= n1500_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9468_q <= n1502_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4073:17  */
  assign n9469_o = clkena_lw ? n9246_o : movem_actiond;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4073:17  */
  always @(posedge clk)
    n9470_q <= n9469_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4073:17  */
  assign n9471_o = {n9380_o, n9406_o, n9403_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9473_q <= n759_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9474_q <= n761_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9475_q <= n1504_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9476_q <= n1506_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9477_q <= n1508_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3239:17  */
  always @(posedge clk)
    n9478_q <= n7945_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9479_q <= n1509_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9480_q <= n1847_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9481_q <= n1511_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9482_q <= n762_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9483_q <= n1513_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:870:17  */
  assign n9484_o = clkena_lw ? n874_o : trap_vector;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:870:17  */
  always @(posedge clk)
    n9485_q <= n9484_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  assign n9486_o = n287_o ? reg_qa : usp;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9487_q <= n9486_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9488_q <= n1514_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9489_q <= n1515_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9490_q <= n1517_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9491_q <= n1849_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9492_q <= n1851_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9493_q <= n1519_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9494_q <= n764_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:743:9  */
  assign n9495_o = {n150_o, n153_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:484:17  */
  assign n9496_o = n157_o ? n162_o : bf_ext_in;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9497_q <= n9496_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9498_q <= n1521_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9499_q <= n1522_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9500_q <= n1523_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9501_q <= n1524_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1254:17  */
  always @(posedge clk)
    n9502_q <= n1578_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9503_q <= n209_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9504_q <= n210_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:484:17  */
  assign n9505_o = {n1705_o, n1702_o, n1708_o};
  assign n9506_o = {1'b0, n1652_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9507_q <= n1525_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9508_q <= n1526_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  assign n9509_o = {1'b0, n1665_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9510_q <= n1527_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9511_q <= n1528_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9512_q <= n9108_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9513_q <= n9110_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9514_q <= n9111_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4008:9  */
  always @(posedge clk)
    n9515_q <= n9112_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:4008:9  */
  assign n9516_o = {n9017_o, n9015_o, n9013_o, n9012_o, n9011_o, n9010_o, n9009_o, n7750_o, n7707_o, n9008_o, n9024_o, n7705_o, n9006_o, n9005_o, n7700_o, n9004_o, n9003_o, n9002_o, n9001_o, n9023_o, n8999_o, n9022_o, n8997_o, n7693_o, n9020_o, n8996_o, n8994_o, n8992_o, n8991_o, n7682_o, n7679_o, n7676_o, n8990_o, n8989_o, n7668_o, n8988_o, n8987_o, n8986_o, n7653_o, n7651_o, n7648_o, n1961_o, n8985_o, n8984_o, n8983_o, n8982_o, n7638_o, n8981_o, n8980_o, n7725_o, n7634_o, n9018_o, n8979_o, n8977_o, n8976_o, n8975_o, n7720_o, n8974_o, n8973_o, n8972_o, n7626_o, n7718_o, n8971_o};
  assign n9517_o = {n7821_o, n7858_o, n7819_o, n7857_o, n7817_o, n7815_o, n7854_o, n7813_o, n7852_o, n7934_o, n7809_o, n7807_o, n7805_o, n7847_o, n7933_o, n7845_o, n7932_o, n9028_o, n9027_o, n9029_o, n7799_o, n7841_o, n7797_o, n7795_o, n7793_o, n7791_o, n7789_o, n7787_o, n7785_o, n7833_o, n7783_o, n7780_o, n7776_o, n7772_o, n7769_o, n7766_o, n7762_o, n7759_o, n7756_o};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1254:17  */
  assign n9518_o = clkena_lw ? n1622_o : exec;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1254:17  */
  always @(posedge clk)
    n9519_q <= n9518_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:3239:17  */
  always @(posedge clk)
    n9520_q <= n7947_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1364:17  */
  always @(posedge clk)
    n9521_q <= n1843_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  always @(posedge clk)
    n9522_q <= n1471_o;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:1053:17  */
  assign n9523_o = {n9521_q, n9522_q};
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:558:35  */
  reg [31:0] regfile[15:0] ; // memory
  initial begin
    regfile[15] = 32'b00000000000000000000000000000000;
    regfile[14] = 32'b00000000000000000000000000000000;
    regfile[13] = 32'b00000000000000000000000000000000;
    regfile[12] = 32'b00000000000000000000000000000000;
    regfile[11] = 32'b00000000000000000000000000000000;
    regfile[10] = 32'b00000000000000000000000000000000;
    regfile[9] = 32'b00000000000000000000000000000000;
    regfile[8] = 32'b00000000000000000000000000000000;
    regfile[7] = 32'b00000000000000000000000000000000;
    regfile[6] = 32'b00000000000000000000000000000000;
    regfile[5] = 32'b00000000000000000000000000000000;
    regfile[4] = 32'b00000000000000000000000000000000;
    regfile[3] = 32'b00000000000000000000000000000000;
    regfile[2] = 32'b00000000000000000000000000000000;
    regfile[1] = 32'b00000000000000000000000000000000;
    regfile[0] = 32'b00000000000000000000000000000000;
    end
  assign n9525_data = regfile[rdindex_b];
  assign n9526_data = regfile[rdindex_a];
  always @(posedge clk)
    if (n283_o)
      regfile[rdindex_a] <= regin;
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:559:35  */
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:558:35  */
  /* ../TG68K.C/TG68KdotC_Kernel.vhd:567:49  */
endmodule

